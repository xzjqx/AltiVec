library verilog;
use verilog.vl_types.all;
entity p405s_mmu_control is
    port(
        MMU_isStatus    : out    vl_logic_vector(0 to 1);
        MMU_isXltValid  : out    vl_logic;
        MMU_icuDsAbort  : out    vl_logic;
        MMU_isRA        : out    vl_logic_vector(22 to 29);
        msrIrL2forITLB  : out    vl_logic;
        LoadRealRaAttr  : out    vl_logic;
        MMU_dsStatus    : out    vl_logic_vector(0 to 7);
        MMU_dcuXltValid : out    vl_logic;
        MMU_dcuUTLBAbort: out    vl_logic;
        MMU_dcuShadowAbort: out    vl_logic;
        MMU_dsRA        : out    vl_logic_vector(22 to 29);
        MMU_wbHold      : out    vl_logic;
        MMU_tlbSXHit    : out    vl_logic;
        MMU_dsStateBorC : out    vl_logic;
        msrDrL2forDTLB  : out    vl_logic;
        MMU_icuIsAbort  : out    vl_logic;
        marRPN          : out    vl_logic_vector(0 to 21);
        marDSize        : out    vl_logic_vector(0 to 6);
        marE            : out    vl_logic;
        marU0           : out    vl_logic;
        marWR           : out    vl_logic;
        marW            : out    vl_logic;
        marG            : out    vl_logic;
        marCacheable    : out    vl_logic;
        marZonePR       : out    vl_logic_vector(0 to 1);
        sprRegE2        : out    vl_logic;
        iccrE1          : out    vl_logic;
        dccrE1          : out    vl_logic;
        sgrE1           : out    vl_logic;
        slerE1          : out    vl_logic;
        skrE1           : out    vl_logic;
        pidE1           : out    vl_logic;
        pidE2           : out    vl_logic;
        zoneE1          : out    vl_logic;
        dcwrE1          : out    vl_logic;
        seldccr         : out    vl_logic;
        seliccr         : out    vl_logic;
        selzone         : out    vl_logic;
        selpid          : out    vl_logic;
        selsgr          : out    vl_logic;
        dearE1          : out    vl_logic;
        dearE2          : out    vl_logic;
        seldcwr         : out    vl_logic;
        selsler         : out    vl_logic;
        selskr          : out    vl_logic;
        seldear         : out    vl_logic;
        MMU_BMCO        : out    vl_logic;
        pidIn_N         : out    vl_logic_vector(0 to 7);
        size_out        : out    vl_logic_vector(0 to 2);
        sprMuxSel       : out    vl_logic_vector(0 to 1);
        wbStorageOp     : in     vl_logic;
        bypassRPN       : out    vl_logic_vector(0 to 21);
        dsStateAfromLatch: out    vl_logic;
        dsStateD        : out    vl_logic;
        dsAddrL2        : out    vl_logic_vector(0 to 2);
        dsrdNotWrt      : out    vl_logic;
        dsEAL           : out    vl_logic_vector(0 to 31);
        dsInvalidate    : out    vl_logic;
        isAddrL2        : out    vl_logic_vector(0 to 1);
        isInvalidate    : out    vl_logic;
        isrdNotWrt      : out    vl_logic;
        isEAL           : out    vl_logic_vector(0 to 21);
        CompE2          : out    vl_logic;
        tlbAddr         : out    vl_logic_vector(0 to 5);
        tagEn           : out    vl_logic;
        dataEn          : out    vl_logic;
        rdWrb           : out    vl_logic;
        indexLookupb    : out    vl_logic;
        EN_ARRAYL1      : out    vl_logic;
        TestComp        : out    vl_logic;
        EN_C1           : out    vl_logic;
        tlb_invalidate  : out    vl_logic;
        tlbE            : out    vl_logic;
        tlbU0           : out    vl_logic;
        DT              : out    vl_logic;
        TID             : out    vl_logic_vector(0 to 7);
        EPN_EA          : out    vl_logic_vector(0 to 21);
        DSIZE           : out    vl_logic_vector(0 to 6);
        RPN             : out    vl_logic_vector(0 to 21);
        tlbV            : out    vl_logic;
        EX              : out    vl_logic;
        WR              : out    vl_logic;
        ZSEL            : out    vl_logic_vector(0 to 3);
        tlbW            : out    vl_logic;
        tlbCacheInhibit : out    vl_logic;
        tlbM            : out    vl_logic;
        tlbG            : out    vl_logic;
        isIReal_N       : out    vl_logic;
        isDsIReal_N     : out    vl_logic;
        isEReal_N       : out    vl_logic;
        isU0Real_N      : out    vl_logic;
        dsIReal_N       : out    vl_logic;
        dsGReal_N       : out    vl_logic;
        dsEReal_N       : out    vl_logic;
        dsU0Real_N      : out    vl_logic;
        wtReqReal_N     : out    vl_logic;
        fetchReq        : in     vl_logic;
        isEA_NEG        : in     vl_logic_vector(0 to 29);
        nonSpecAcc      : in     vl_logic;
        isAbort         : in     vl_logic;
        cntxSync        : in     vl_logic;
        msrIR           : in     vl_logic;
        isNP            : in     vl_logic;
        isCA            : in     vl_logic;
        EoOdd           : in     vl_logic;
        CancelData      : in     vl_logic;
        icuOp           : in     vl_logic;
        isNewLine       : in     vl_logic;
        msrPR           : in     vl_logic;
        msrDR           : in     vl_logic;
        LdNotSt         : in     vl_logic;
        wbAbort         : in     vl_logic;
        dcuOp           : in     vl_logic;
        dsMmuOp         : in     vl_logic_vector(0 to 3);
        dsEA_N          : in     vl_logic_vector(0 to 31);
        ICU_dsCA        : in     vl_logic;
        DCU_CA          : in     vl_logic;
        cdbcrFDK        : in     vl_logic;
        dcuLoad         : in     vl_logic;
        dcuStore        : in     vl_logic;
        dcbz            : in     vl_logic;
        dcba            : in     vl_logic;
        VCT_mmuExeSuppress: in     vl_logic;
        IFB_exeFlush    : in     vl_logic;
        PCL_mmuExeAbort : in     vl_logic;
        tlbSX           : in     vl_logic;
        tlbWE           : in     vl_logic;
        tlbRE           : in     vl_logic;
        tlbWC           : in     vl_logic;
        exeTlbOp        : in     vl_logic;
        sprAddr         : in     vl_logic_vector(4 to 9);
        SprDcd          : in     vl_logic_vector(0 to 8);
        sprData         : in     vl_logic_vector(0 to 31);
        mtSPR           : in     vl_logic;
        mfSPR           : in     vl_logic;
        sprHold         : in     vl_logic;
        VCT_dearE2      : in     vl_logic;
        iccrL2          : in     vl_logic_vector(0 to 31);
        dccrL2          : in     vl_logic_vector(0 to 31);
        dcwrL2          : in     vl_logic_vector(0 to 31);
        slerL2          : in     vl_logic_vector(0 to 31);
        skrL2           : in     vl_logic_vector(0 to 31);
        sgrL2           : in     vl_logic_vector(0 to 31);
        pidL2           : in     vl_logic_vector(0 to 7);
        zoneL2          : in     vl_logic_vector(0 to 31);
        UTLB_DSize      : in     vl_logic_vector(0 to 6);
        UTLB_EPN        : in     vl_logic_vector(0 to 21);
        UTLB_V          : in     vl_logic;
        UTLB_E          : in     vl_logic;
        UTLB_U0         : in     vl_logic;
        UTLB_TID        : in     vl_logic_vector(0 to 7);
        UTLB_Miss       : in     vl_logic;
        UTLB_RPN        : in     vl_logic_vector(0 to 21);
        UTLB_EX         : in     vl_logic;
        UTLB_WR         : in     vl_logic;
        UTLB_ZSEL       : in     vl_logic_vector(0 to 3);
        UTLB_W          : in     vl_logic;
        UTLB_CacheInhibit: in     vl_logic;
        UTLB_G          : in     vl_logic;
        dtlbMiss        : in     vl_logic;
        DTLB_zonePR     : in     vl_logic_vector(0 to 1);
        DTLB_WR         : in     vl_logic;
        DTLB_U0         : in     vl_logic;
        DTLB_I          : in     vl_logic;
        DTLB_W          : in     vl_logic;
        itlbMiss        : in     vl_logic;
        PCL_wbHoldnonErr: in     vl_logic;
        exeStorageOp    : in     vl_logic;
        resetL2         : in     vl_logic;
        CB              : in     vl_logic;
        TestM1          : in     vl_logic;
        TestM3          : in     vl_logic;
        LSSD_ArrayCClk_buf: in     vl_logic;
        BIST_wrEn       : in     vl_logic;
        BIST_rdEn       : in     vl_logic;
        BIST_addr       : in     vl_logic_vector(0 to 5);
        BIST_lookupEn   : in     vl_logic;
        BIST_epn_ea     : in     vl_logic_vector(0 to 21);
        BIST_DSize      : in     vl_logic_vector(0 to 6);
        BIST_TID        : in     vl_logic_vector(0 to 7);
        BIST_data       : in     vl_logic_vector(0 to 1);
        BIST_DT         : in     vl_logic;
        BIST_V          : in     vl_logic;
        BIST_invalidate : in     vl_logic;
        ABIST_test      : in     vl_logic;
        EN_ARRAYL1_preTestM3: out    vl_logic;
        UTLB_DT         : in     vl_logic;
        MMU_tlbREParityErr: out    vl_logic;
        MMU_tlbSXParityErr: out    vl_logic;
        MMU_dsParityErr : out    vl_logic;
        MMU_isParityErr : out    vl_logic;
        tagPar1         : out    vl_logic;
        tagPar2         : out    vl_logic;
        tagPar3         : out    vl_logic;
        tagPar4         : out    vl_logic;
        ramPar1         : out    vl_logic;
        ramPar2         : out    vl_logic;
        UTLB_T1         : in     vl_logic;
        UTLB_T2         : in     vl_logic;
        UTLB_T3         : in     vl_logic;
        UTLB_T4         : in     vl_logic;
        UTLB_R1         : in     vl_logic;
        UTLB_R2         : in     vl_logic;
        UTLB_M          : in     vl_logic;
        ICU_CCR1TLBE    : in     vl_logic;
        ICU_CCR0TPE     : in     vl_logic
    );
end p405s_mmu_control;
