library verilog;
use verilog.vl_types.all;
entity p405s_brEquations is
    port(
        pfb0Branch      : out    vl_logic;
        nxtPfb0FirstCycle: out    vl_logic;
        pfb0Bc          : out    vl_logic;
        pfb0Target_Neg  : out    vl_logic;
        pfb0PredictionHolding: out    vl_logic;
        nxtDcdPfb0Prediction: out    vl_logic;
        dcdPredict      : out    vl_logic;
        dcdPrediction   : out    vl_logic;
        nxtExeDcdPrediction_Neg: out    vl_logic;
        dcdCorrect_Neg  : out    vl_logic;
        dcdCtrEq0       : out    vl_logic;
        nxtDcdFirstCycle: out    vl_logic;
        dcdHold_Neg     : out    vl_logic;
        dcdPredictHolding: out    vl_logic;
        nxtExeDcdPredict: out    vl_logic;
        dcdPredictionHolding: out    vl_logic;
        exeCorrect      : out    vl_logic;
        exeCorrect_Neg  : out    vl_logic;
        exeBrAndLink    : out    vl_logic;
        nxtExeFirstCycle: out    vl_logic;
        exeCrtBpntLrCtr : out    vl_logic;
        branchTarCrt    : out    vl_logic;
        IFB_exeDbgBrTaken: out    vl_logic;
        dcdCrtE2        : out    vl_logic;
        dcdCrtMuxSel    : out    vl_logic;
        exeCrtE2        : out    vl_logic;
        exeCrtMuxSel    : out    vl_logic_vector(0 to 1);
        pfb0PlaB        : in     vl_logic;
        pfb0PlaBc       : in     vl_logic;
        pfb0PriOp_5     : in     vl_logic;
        pfb0SecOp_0     : in     vl_logic;
        pfb0DataBO_0    : in     vl_logic;
        pfb0DataBO_2    : in     vl_logic;
        pfb0DataBO_4    : in     vl_logic;
        pfb0DataBD_0    : in     vl_logic;
        pfb0FullL2      : in     vl_logic;
        pfb0FirstCycleL2: in     vl_logic;
        pfb0PredictionHoldingL2: in     vl_logic;
        dcdPlaB         : in     vl_logic;
        dcdPlaBc        : in     vl_logic;
        dcdPlaMtspr     : in     vl_logic;
        dcdDataBO_0     : in     vl_logic;
        dcdDataBO_2     : in     vl_logic;
        dcdDataBO_4     : in     vl_logic;
        dcdDataBD_0     : in     vl_logic;
        dcdDataL2       : in     vl_logic_vector(11 to 20);
        dcdPriOp_5      : in     vl_logic;
        dcdSecOp_0      : in     vl_logic;
        dcdDataLK       : in     vl_logic;
        dcdPfb0PredictionL2: in     vl_logic;
        dcdPfb0BranchL2 : in     vl_logic;
        dcdPfb0BcL2     : in     vl_logic;
        dcdCrtBpntLrCtr : out    vl_logic;
        dcdCondOK       : in     vl_logic;
        dcdTarget_Neg   : in     vl_logic;
        dcdFullL2       : in     vl_logic;
        dcdFirstCycleL2 : in     vl_logic;
        dcdClear        : in     vl_logic;
        dcdFlush        : in     vl_logic;
        dcdPredictHoldingL2: in     vl_logic;
        dcdPredictionHoldingL2: in     vl_logic;
        exeBL2          : in     vl_logic;
        exeBcL2         : in     vl_logic;
        exeMtCtrL2      : in     vl_logic;
        exeDataBO_2     : in     vl_logic;
        exeDataLKL2     : in     vl_logic;
        exeFullL2       : in     vl_logic;
        exeFirstCycleL2 : in     vl_logic;
        exeDcdPredictL2 : in     vl_logic;
        exeDcdPrediction_NegL2: in     vl_logic;
        exeCondOK_Neg   : in     vl_logic;
        exe2Cr0EnL2     : in     vl_logic;
        exeCrUpdateL2   : in     vl_logic;
        exeCtrUpForBcctrL2: in     vl_logic;
        exeLrUpdateL2   : in     vl_logic;
        exeDataBr_5L2   : in     vl_logic;
        ctrEq1L2        : in     vl_logic;
        ctrEq2L2        : in     vl_logic;
        PCL_dcdHoldForIFB: in     vl_logic;
        PCL_exeIarHold  : in     vl_logic;
        tracePipeHold   : in     vl_logic
    );
end p405s_brEquations;
