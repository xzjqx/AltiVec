library verilog;
use verilog.vl_types.all;
entity p405s_MMU_top is
    port(
        CAR_U0Attr      : out    vl_logic;
        CAR_cacheable   : out    vl_logic;
        CAR_endian      : out    vl_logic;
        CAR_guarded     : out    vl_logic;
        CAR_writethru   : out    vl_logic;
        MMU_BMCO        : out    vl_logic;
        MMU_apuWbEndian : out    vl_logic;
        MMU_dcuShadowAbort: out    vl_logic;
        MMU_dcuUTLBAbort: out    vl_logic;
        MMU_dcuXltValid : out    vl_logic;
        MMU_diagOut     : out    vl_logic_vector(0 to 2);
        MMU_dsRA        : out    vl_logic_vector(0 to 29);
        MMU_dsStateBorC : out    vl_logic;
        MMU_dsStatus    : out    vl_logic_vector(0 to 7);
        MMU_dsocmABus   : out    vl_logic_vector(0 to 29);
        MMU_dsocmCacheable: out    vl_logic;
        MMU_dsocmGuarded: out    vl_logic;
        MMU_dsocmU0Attr : out    vl_logic;
        MMU_dsocmXltValid: out    vl_logic;
        MMU_icuDsAbort  : out    vl_logic;
        MMU_icuIsAbort  : out    vl_logic;
        MMU_isCacheable_NEG: out    vl_logic_vector(0 to 2);
        MMU_isDsCacheableL2: out    vl_logic;
        MMU_isDsEndianL2: out    vl_logic;
        MMU_isDsU0AttrL2: out    vl_logic;
        MMU_isDsXltValidL2: out    vl_logic;
        MMU_isEndian    : out    vl_logic;
        MMU_isRA_NEG    : out    vl_logic_vector(0 to 29);
        MMU_isStatus    : out    vl_logic_vector(0 to 1);
        MMU_isU0Attr    : out    vl_logic;
        MMU_isXltValid  : out    vl_logic;
        MMU_isocmCacheable: out    vl_logic;
        MMU_isocmU0Attr : out    vl_logic;
        MMU_isocmXltValid: out    vl_logic;
        MMU_rdarDsRAL2  : out    vl_logic_vector(0 to 29);
        MMU_sprData     : out    vl_logic_vector(0 to 31);
        MMU_tlbSXHit    : out    vl_logic;
        MMU_wbHold      : out    vl_logic;
        CAR_mmuAttr_E1  : in     vl_logic;
        CAR_mmuAttr_E2  : in     vl_logic;
        CB              : in     vl_logic;
        DCU_CA          : in     vl_logic;
        EXE_dsEA_NEG    : in     vl_logic_vector(0 to 31);
        EXE_dsEaCP_NEG  : in     vl_logic_vector(0 to 7);
        EXE_eaARegBuf   : in     vl_logic_vector(0 to 21);
        EXE_eaBRegBuf   : in     vl_logic_vector(0 to 21);
        EXE_mmuIcuSprData: in     vl_logic_vector(0 to 31);
        EXE_sprAddr     : in     vl_logic_vector(4 to 9);
        ICU_CCR0DDK     : in     vl_logic;
        ICU_EoOdd       : in     vl_logic;
        ICU_dsCA        : in     vl_logic;
        ICU_isCA        : in     vl_logic;
        ICU_mmuRdarE2   : in     vl_logic;
        IFB_cntxSync    : in     vl_logic;
        IFB_exeFlush    : in     vl_logic;
        IFB_fetchReq    : in     vl_logic;
        IFB_icuCancelData: in     vl_logic;
        IFB_isAbort     : in     vl_logic;
        IFB_isEA        : in     vl_logic_vector(0 to 29);
        IFB_isNL        : in     vl_logic;
        IFB_isNP        : in     vl_logic;
        IFB_nonSpecAcc  : in     vl_logic;
        LSSD_TestM1     : in     vl_logic;
        LSSD_TestM3     : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        MMU_BIST_Scanin : in     vl_logic;
        MMU_scanIn      : in     vl_logic_vector(0 to 3);
        PCL_dcba        : in     vl_logic;
        PCL_dcbz        : in     vl_logic;
        PCL_dcuLoad     : in     vl_logic;
        PCL_dcuOp       : in     vl_logic;
        PCL_dcuStore    : in     vl_logic;
        PCL_dsMmuOp     : in     vl_logic_vector(0 to 3);
        PCL_exeStorageOp: in     vl_logic;
        PCL_exeTlbOp    : in     vl_logic;
        PCL_icuOp       : in     vl_logic;
        PCL_ldNotSt     : in     vl_logic;
        PCL_mfSPR       : in     vl_logic;
        PCL_mmuExeAbort : in     vl_logic;
        PCL_mmuIcuSprHold: in     vl_logic;
        PCL_mmuSprDcd   : in     vl_logic_vector(0 to 8);
        PCL_mtSPR       : in     vl_logic;
        PCL_tlbRE       : in     vl_logic;
        PCL_tlbSX       : in     vl_logic;
        PCL_tlbWE       : in     vl_logic;
        PCL_tlbWS       : in     vl_logic;
        PCL_wbHoldNonErr: in     vl_logic;
        PCL_wbStorageOp : in     vl_logic;
        VCT_dcuWbAbort  : in     vl_logic;
        VCT_dearE2      : in     vl_logic;
        VCT_mmuExeSuppress: in     vl_logic;
        VCT_msrDR       : in     vl_logic;
        VCT_msrIR       : in     vl_logic;
        VCT_msrPR       : in     vl_logic;
        resetCore       : in     vl_logic;
        testmode        : in     vl_logic;
        MMU_tlbREParityErr: out    vl_logic;
        MMU_tlbSXParityErr: out    vl_logic;
        MMU_dsParityErr : out    vl_logic;
        MMU_isParityErr : out    vl_logic;
        ICU_CCR0PRS     : in     vl_logic;
        BIST_pepsPF     : out    vl_logic_vector(0 to 2);
        ICU_CCR1TLBE    : in     vl_logic;
        ICU_CCR0TPE     : in     vl_logic;
        LSSD_EVS        : in     vl_logic;
        BISTCE0STCLK    : in     vl_logic;
        BISTCE1ENABLE   : in     vl_logic;
        LSSD_BISTCClk   : in     vl_logic;
        BIST_Done       : out    vl_logic;
        resetMemBist    : out    vl_logic
    );
end p405s_MMU_top;
