library verilog;
use verilog.vl_types.all;
entity p405s_adm_top is
    port(
        EXE_admMco      : out    vl_logic;
        EXE_divMco      : out    vl_logic;
        EXE_multMco     : out    vl_logic;
        aRegMuxSel      : out    vl_logic_vector(0 to 1);
        aRegZ4dndSEIn   : out    vl_logic_vector(0 to 4);
        addCA           : out    vl_logic;
        addOV           : out    vl_logic;
        admCcBits       : out    vl_logic_vector(0 to 2);
        admCcMuxSel     : out    vl_logic_vector(0 to 1);
        admOut          : out    vl_logic_vector(0 to 31);
        bRegMuxSel      : out    vl_logic_vector(0 to 1);
        divNxtToLastSt  : out    vl_logic;
        divOV           : out    vl_logic;
        divPathEn       : out    vl_logic;
        macOV           : out    vl_logic;
        macOVSat_NEG    : out    vl_logic;
        macSatValue     : out    vl_logic_vector(0 to 2);
        multHiEOAnsCc   : out    vl_logic_vector(0 to 2);
        multLo4CycAnsCc : out    vl_logic_vector(0 to 2);
        multLo5CycAnsCc : out    vl_logic_vector(0 to 2);
        multOV          : out    vl_logic;
        nxtQ            : out    vl_logic;
        nxtQ_NEG        : out    vl_logic;
        resetL2         : out    vl_logic;
        sRegMuxSel      : out    vl_logic_vector(0 to 1);
        srmMuxSel       : out    vl_logic_vector(0 to 5);
        trap            : out    vl_logic;
        CB              : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        PCL_aPortRregBypass: in     vl_logic;
        PCL_addFour     : in     vl_logic;
        PCL_bPortLitGenSel: in     vl_logic;
        PCL_bPortRregBypass: in     vl_logic;
        PCL_dcdAregLoadUse: in     vl_logic;
        PCL_dcdBregLoadUse: in     vl_logic;
        PCL_dcdHotCIn   : in     vl_logic;
        PCL_dcdMdSelQ   : in     vl_logic;
        PCL_dcdMrSelQ   : in     vl_logic;
        PCL_dcdSregLoadUse: in     vl_logic;
        PCL_dcdSrmBpSel : in     vl_logic_vector(0 to 2);
        PCL_dcdXerCa    : in     vl_logic;
        PCL_exe2AccRegMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exe2Hold    : in     vl_logic;
        PCL_exe2MacEn   : in     vl_logic;
        PCL_exe2MacOrMultEnForMS: in     vl_logic_vector(0 to 1);
        PCL_exe2MacOrMultEn_NEG: in     vl_logic_vector(0 to 1);
        PCL_exe2MacSat  : in     vl_logic;
        PCL_exe2MultEn  : in     vl_logic;
        PCL_exe2MultHiWd: in     vl_logic;
        PCL_exe2NegMac  : in     vl_logic;
        PCL_exe2SignedOp: in     vl_logic;
        PCL_exe2XerOvEn : in     vl_logic;
        PCL_exeAddSgndOp_NEG: in     vl_logic_vector(0 to 1);
        PCL_exeAdmCntl  : in     vl_logic_vector(0 to 3);
        PCL_exeAregLoadUse: in     vl_logic;
        PCL_exeBregLoadUse: in     vl_logic;
        PCL_exeCmplmntA : in     vl_logic;
        PCL_exeCmplmntA_NEG: in     vl_logic;
        PCL_exeDivEn    : in     vl_logic;
        PCL_exeDivEnForLSSD: in     vl_logic;
        PCL_exeDivEnForMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exeDivEn_NEG: in     vl_logic;
        PCL_exeDivSgndOp: in     vl_logic;
        PCL_exeDvcHold  : in     vl_logic;
        PCL_exeLoadUseHold: in     vl_logic;
        PCL_exeMacEn    : in     vl_logic;
        PCL_exeMultEn   : in     vl_logic;
        PCL_exeMultEnForMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exeMultEn_NEG: in     vl_logic_vector(0 to 1);
        PCL_exeNegMac   : in     vl_logic;
        PCL_exeSregLoadUse: in     vl_logic;
        PCL_exeSrmBpSel : in     vl_logic_vector(0 to 2);
        PCL_exeXerOvEn  : in     vl_logic;
        PCL_gateZeroToAreg: in     vl_logic;
        PCL_gateZeroToSreg: in     vl_logic;
        PCL_holdCIn     : in     vl_logic;
        PCL_holdMdMr    : in     vl_logic;
        PCL_sPortRregBypass: in     vl_logic;
        PCL_wbHold      : in     vl_logic;
        aReg_NEG        : in     vl_logic_vector(0 to 31);
        bReg_NEG        : in     vl_logic_vector(0 to 31);
        coreReset       : in     vl_logic;
        deterministicMult: in     vl_logic;
        exeMacOrMultEn_NEG: in     vl_logic;
        nxtXerCa        : in     vl_logic;
        rRegBypassForAccReg: in     vl_logic_vector(0 to 31);
        sBus            : in     vl_logic_vector(0 to 31);
        trapCond        : in     vl_logic_vector(0 to 4);
        PCL_exeDvcOrParityHold: in     vl_logic
    );
end p405s_adm_top;
