library verilog;
use verilog.vl_types.all;
entity p405s_jtg_top is
    port(
        JTG_TDO         : out    vl_logic;
        JTG_captureDR   : out    vl_logic;
        JTG_dbdrPulse   : out    vl_logic;
        JTG_dbgWaitEn   : out    vl_logic;
        JTG_extest      : out    vl_logic;
        JTG_freezeTimers: out    vl_logic;
        JTG_iCacheWr_NEG: out    vl_logic;
        JTG_inst        : out    vl_logic_vector(0 to 31);
        JTG_instBuf     : out    vl_logic_vector(0 to 31);
        JTG_pgmOut      : out    vl_logic;
        JTG_resetChipReq: out    vl_logic;
        JTG_resetCoreReq: out    vl_logic;
        JTG_resetDBSR   : out    vl_logic;
        JTG_resetSystemReq: out    vl_logic;
        JTG_shiftDR     : out    vl_logic;
        JTG_sprDataBus  : out    vl_logic_vector(0 to 31);
        JTG_step        : out    vl_logic;
        JTG_stepUPD     : out    vl_logic;
        JTG_stopReq     : out    vl_logic;
        JTG_stuff       : out    vl_logic;
        JTG_stuffUPD    : out    vl_logic;
        JTG_tDOEnable   : out    vl_logic;
        JTG_uncondEvent : out    vl_logic;
        JTG_updateDR    : out    vl_logic;
        CB              : in     vl_logic;
        CPM_coreClkOff  : in     vl_logic;
        DBG_DE          : in     vl_logic;
        DBG_UDE         : in     vl_logic;
        DBG_resetChip   : in     vl_logic;
        DBG_resetCore   : in     vl_logic;
        DBG_resetSystem : in     vl_logic;
        EXE_sprDataBus  : in     vl_logic_vector(0 to 31);
        ICU_sleepReq    : in     vl_logic;
        IFB_msrWE       : in     vl_logic;
        IFB_rstStepPend : in     vl_logic;
        IFB_rstStuffPend: in     vl_logic;
        IFB_stopAck     : in     vl_logic;
        JTGEX_BndScanTDO: in     vl_logic;
        JTGEX_TCK       : in     vl_logic;
        JTGEX_TDI       : in     vl_logic;
        JTGEX_TMS       : in     vl_logic;
        JTGEX_TRST_NEG  : in     vl_logic;
        PCL_exeMfspr    : in     vl_logic;
        PCL_exeMtspr    : in     vl_logic;
        PCL_exeSprHold  : in     vl_logic;
        PCL_jtgSprDcd   : in     vl_logic;
        PLB_jtgHoldAck  : in     vl_logic;
        TIM_wdChipRst   : in     vl_logic;
        TIM_wdCoreRst   : in     vl_logic;
        TIM_wdSysRst    : in     vl_logic;
        VCT_msrDWE      : in     vl_logic;
        VCT_srr1DWE     : in     vl_logic;
        VCT_srr3DWE     : in     vl_logic;
        VCT_stuffStepSup: in     vl_logic;
        VCT_sxr         : in     vl_logic_vector(0 to 11);
        XXX_coreReset   : in     vl_logic;
        XXX_jtgHalt     : in     vl_logic;
        XXX_systemReset : in     vl_logic;
        jtgDiagBus1     : in     vl_logic_vector(0 to 31);
        jtgDiagBus2     : in     vl_logic_vector(0 to 31);
        jtgDiagBus3     : in     vl_logic_vector(0 to 31)
    );
end p405s_jtg_top;
