library verilog;
use verilog.vl_types.all;
entity p405s_branchCntl is
    port(
        IFB_exeCorrect  : out    vl_logic;
        IFB_exeDbgBrTaken: out    vl_logic;
        branchTarCrt    : out    vl_logic;
        dcdCorrect_Neg  : out    vl_logic;
        dcdCrtBpntLrCtr : out    vl_logic;
        dcdCrtE2        : out    vl_logic;
        dcdCrtMuxSel    : out    vl_logic;
        dcdTarget_Neg   : out    vl_logic;
        exeBrAndLink    : out    vl_logic;
        exeCorrect_Neg  : out    vl_logic;
        exeCrtBpntLrCtr : out    vl_logic;
        exeCrtE2        : out    vl_logic;
        exeCrtMuxSel    : out    vl_logic_vector(0 to 1);
        pfb0Target_Neg  : out    vl_logic;
        CB              : in     vl_logic;
        PCL_dcdHoldForIFB: in     vl_logic;
        PCL_exeIarHold  : in     vl_logic;
        crL2            : in     vl_logic_vector(0 to 31);
        ctrEq1L2        : in     vl_logic;
        ctrEq2L2        : in     vl_logic;
        dcdClear        : in     vl_logic;
        dcdDataBD_0     : in     vl_logic;
        dcdDataBI       : in     vl_logic_vector(0 to 4);
        dcdDataBO       : in     vl_logic_vector(0 to 4);
        dcdDataL2       : in     vl_logic_vector(11 to 20);
        dcdDataLK       : in     vl_logic;
        dcdFlush        : in     vl_logic;
        dcdFullL2       : in     vl_logic;
        dcdPlaB         : in     vl_logic;
        dcdPlaBc        : in     vl_logic;
        dcdPlaMtspr     : in     vl_logic;
        dcdPriOp_5      : in     vl_logic;
        dcdSecOp_0      : in     vl_logic;
        exe2Cr0EnL2     : in     vl_logic;
        exeBL2          : in     vl_logic;
        exeBcL2         : in     vl_logic;
        exeCrUpdateL2   : in     vl_logic;
        exeCtrUpForBcctrL2: in     vl_logic;
        exeDataBrBIL2   : in     vl_logic_vector(0 to 4);
        exeDataBrBOL2   : in     vl_logic_vector(0 to 3);
        exeDataBr_5L2   : in     vl_logic;
        exeDataLKL2     : in     vl_logic;
        exeFullL2       : in     vl_logic;
        exeLrUpdateL2   : in     vl_logic;
        exeMtCtrL2      : in     vl_logic;
        pfb0DataBD_0    : in     vl_logic;
        pfb0DataBO_0    : in     vl_logic;
        pfb0DataBO_2    : in     vl_logic;
        pfb0DataBO_4    : in     vl_logic;
        pfb0FullL2      : in     vl_logic;
        pfb0PlaB        : in     vl_logic;
        pfb0PlaBc       : in     vl_logic;
        pfb0PriOp_5     : in     vl_logic;
        pfb0SecOp_0     : in     vl_logic;
        tracePipeHold   : in     vl_logic
    );
end p405s_branchCntl;
