library verilog;
use verilog.vl_types.all;
entity top_class_based is
end top_class_based;
