library verilog;
use verilog.vl_types.all;
entity p405s_cpu_top is
    port(
        C405_jtgCaptureDR: out    vl_logic;
        C405_jtgExtest  : out    vl_logic;
        C405_jtgPlbDcuPriorityAdjust: out    vl_logic;
        C405_jtgShiftDR : out    vl_logic;
        C405_jtgTDO     : out    vl_logic;
        C405_jtgTDOEn   : out    vl_logic;
        C405_jtgUpdateDR: out    vl_logic;
        C405_rstChipResetReq: out    vl_logic;
        C405_rstCoreResetReq: out    vl_logic;
        C405_rstSystemResetReq: out    vl_logic;
        CPU_TEType      : out    vl_logic_vector(0 to 10);
        Core_lssdScanOut: out    vl_logic_vector(10 to 31);
        DCU_parityError : in     vl_logic;
        DCU_FlushParityError: in     vl_logic;
        EXE_apuLoadData : out    vl_logic_vector(0 to 31);
        EXE_dcrAddr     : out    vl_logic_vector(0 to 9);
        EXE_dcrDataBus  : out    vl_logic_vector(0 to 31);
        EXE_dcuData     : out    vl_logic_vector(0 to 31);
        EXE_dsEA_NEG    : out    vl_logic_vector(0 to 31);
        EXE_dsEaCP      : out    vl_logic_vector(0 to 7);
        EXE_eaARegBuf   : out    vl_logic_vector(0 to 21);
        EXE_eaBRegBuf   : out    vl_logic_vector(0 to 21);
        EXE_icuSprDcds  : out    vl_logic_vector(0 to 2);
        EXE_mmuIcuSprDataBus: out    vl_logic_vector(0 to 31);
        EXE_raData      : out    vl_logic_vector(0 to 31);
        EXE_rbData      : out    vl_logic_vector(0 to 31);
        ICU_parityErrE  : in     vl_logic;
        ICU_parityErrO  : in     vl_logic;
        ICU_tagParityErr: in     vl_logic;
        ICU_CCR0DPP     : in     vl_logic;
        ICU_CCR0DPE     : in     vl_logic;
        ICU_CCR0IPE     : in     vl_logic;
        ICU_CCR0TPE     : in     vl_logic;
        EXE_sprAddr     : out    vl_logic_vector(4 to 9);
        EXE_xerCa       : out    vl_logic;
        IFB_TE          : out    vl_logic;
        IFB_cntxSync    : out    vl_logic;
        IFB_cntxSyncOCM : out    vl_logic;
        IFB_coreSleepReq: out    vl_logic;
        IFB_dcdFullApuL2: out    vl_logic;
        IFB_exeFlush    : out    vl_logic;
        IFB_extStopAck  : out    vl_logic;
        IFB_fetchReq    : out    vl_logic;
        IFB_icuCancelDataL2: out    vl_logic;
        IFB_isAbortForICU: out    vl_logic_vector(0 to 2);
        IFB_isAbortForMMU: out    vl_logic;
        IFB_isEA        : out    vl_logic_vector(0 to 29);
        IFB_isNL        : out    vl_logic;
        IFB_isNP        : out    vl_logic;
        IFB_isOcmAbus_Neg: out    vl_logic_vector(0 to 29);
        IFB_nonSpecAcc  : out    vl_logic;
        IFB_ocmAbort    : out    vl_logic;
        IFB_regDcdApuL2 : out    vl_logic_vector(0 to 31);
        IFB_wbIar       : out    vl_logic_vector(0 to 29);
        JTG_iCacheWr    : out    vl_logic;
        JTG_instBuf     : out    vl_logic_vector(0 to 31);
        MMU_tlbREParityErr: in     vl_logic;
        MMU_tlbSXParityErr: in     vl_logic;
        MMU_dsParityErr : in     vl_logic;
        MMU_isParityErr : in     vl_logic;
        PCL_apuExeWdCnt : out    vl_logic_vector(0 to 1);
        PCL_apuLoadDV   : out    vl_logic;
        PCL_apuWbHold   : out    vl_logic;
        PCL_dcdHoldForApu: out    vl_logic;
        PCL_dcuByteEn   : out    vl_logic_vector(0 to 3);
        PCL_dcuOp       : out    vl_logic_vector(0 to 11);
        PCL_dcuOp_early : out    vl_logic_vector(0 to 2);
        PCL_dsMmuOp     : out    vl_logic_vector(0 to 3);
        PCL_dsOcmByteEn : out    vl_logic_vector(0 to 3);
        PCL_exeAbort    : out    vl_logic;
        PCL_exeFlushForApu: out    vl_logic;
        PCL_exeHoldForApu: out    vl_logic;
        PCL_exeLdNotSt  : out    vl_logic;
        PCL_exeStorageOp: out    vl_logic;
        PCL_exeStringMultiple: out    vl_logic;
        PCL_exeTlbOp    : out    vl_logic;
        PCL_icuOp       : out    vl_logic_vector(0 to 3);
        PCL_mfDCR       : out    vl_logic;
        PCL_mfSPR       : out    vl_logic;
        PCL_mmuExeAbort : out    vl_logic;
        PCL_mmuIcuSprHold: out    vl_logic;
        PCL_mmuSprDcd   : out    vl_logic_vector(0 to 8);
        PCL_mtDCR       : out    vl_logic;
        PCL_mtSPR       : out    vl_logic;
        PCL_ocmAbortReq : out    vl_logic;
        PCL_stSteerCntl : out    vl_logic_vector(0 to 9);
        PCL_tlbRE       : out    vl_logic;
        PCL_tlbSX       : out    vl_logic;
        PCL_tlbWE       : out    vl_logic;
        PCL_tlbWS       : out    vl_logic;
        PCL_trcLoadDV   : out    vl_logic;
        PCL_wbComplete  : out    vl_logic;
        PCL_wbFull      : out    vl_logic;
        PCL_wbHoldNonErr: out    vl_logic;
        PCL_wbStorageOp : out    vl_logic;
        TIM_timerResetL2: out    vl_logic;
        TRC_evenESBusL2 : out    vl_logic_vector(0 to 1);
        TRC_oddCycle    : out    vl_logic;
        TRC_oddESBusL2  : out    vl_logic_vector(0 to 1);
        TRC_tsBusL2     : out    vl_logic_vector(0 to 3);
        VCT_apuWbFlush  : out    vl_logic;
        VCT_dcuWbAbort  : out    vl_logic;
        VCT_dearE2      : out    vl_logic;
        VCT_errorOut    : out    vl_logic;
        VCT_icuWbAbort  : out    vl_logic;
        VCT_mmuExeSuppress: out    vl_logic;
        VCT_mmuWbAbort  : out    vl_logic;
        VCT_msrCE       : out    vl_logic;
        VCT_msrDR       : out    vl_logic;
        VCT_msrEE       : out    vl_logic;
        VCT_msrFE0      : out    vl_logic;
        VCT_msrFE1      : out    vl_logic;
        VCT_msrIR       : out    vl_logic;
        VCT_msrPR       : out    vl_logic;
        VCT_msrWE       : out    vl_logic;
        VCT_timerIntrp  : out    vl_logic;
        APU_dcdApuOp    : in     vl_logic;
        APU_dcdExeLdDepend: in     vl_logic;
        APU_dcdForceAlgn: in     vl_logic;
        APU_dcdForceBESteering: in     vl_logic;
        APU_dcdFpuOp    : in     vl_logic;
        APU_dcdGprWr    : in     vl_logic;
        APU_dcdLdStByte : in     vl_logic;
        APU_dcdLdStDw   : in     vl_logic;
        APU_dcdLdStHw   : in     vl_logic;
        APU_dcdLdStQw   : in     vl_logic;
        APU_dcdLdStWd   : in     vl_logic;
        APU_dcdLoad     : in     vl_logic;
        APU_dcdLwbLdDepend: in     vl_logic;
        APU_dcdPrivOp   : in     vl_logic;
        APU_dcdRaEn     : in     vl_logic;
        APU_dcdRbEn     : in     vl_logic;
        APU_dcdRc       : in     vl_logic;
        APU_dcdStore    : in     vl_logic;
        APU_dcdTrapBE   : in     vl_logic;
        APU_dcdTrapLE   : in     vl_logic;
        APU_dcdUpdate   : in     vl_logic;
        APU_dcdValidOp  : in     vl_logic;
        APU_dcdWbLdDepend: in     vl_logic;
        APU_dcdXerCAEn  : in     vl_logic;
        APU_dcdXerOVEn  : in     vl_logic;
        APU_exception   : in     vl_logic;
        APU_exeBlkingMco: in     vl_logic;
        APU_exeBusy     : in     vl_logic;
        APU_exeCa       : in     vl_logic;
        APU_exeCr       : in     vl_logic_vector(0 to 3);
        APU_exeCrField  : in     vl_logic_vector(0 to 2);
        APU_exeNonBlkingMco: in     vl_logic;
        APU_exeOv       : in     vl_logic;
        APU_exeResult   : in     vl_logic_vector(0 to 31);
        APU_sleepReq    : in     vl_logic;
        C405_timerTick  : in     vl_logic;
        CAR_cacheable   : in     vl_logic;
        CAR_endian      : in     vl_logic;
        CB              : in     vl_logic;
        TimerClk        : in     vl_logic;
        CPM_coreClkOff  : in     vl_logic;
        DBG_c405DebugHalt: in     vl_logic;
        DBG_c405ExtBusHoldAck: in     vl_logic;
        DCU_CA          : in     vl_logic;
        DCU_DA          : in     vl_logic;
        DCU_SCL2        : in     vl_logic;
        DCU_SDQ_mod     : in     vl_logic_vector(0 to 31);
        DCU_carByteEn   : in     vl_logic_vector(0 to 3);
        DCU_data_NEG    : in     vl_logic_vector(0 to 31);
        DCU_diagBus     : in     vl_logic_vector(0 to 20);
        DCU_firstCycCarStXltV: in     vl_logic;
        DCU_pclOcmWait  : in     vl_logic;
        DCU_sleepReq    : in     vl_logic;
        EIC_critIntrp   : in     vl_logic;
        EIC_extIntrp    : in     vl_logic;
        FPU_exception   : in     vl_logic;
        ICU_EO          : in     vl_logic_vector(0 to 1);
        ICU_GPRC        : in     vl_logic;
        ICU_LDBE        : in     vl_logic;
        ICU_diagBus     : in     vl_logic_vector(0 to 22);
        ICU_dsCA        : in     vl_logic;
        ICU_ifbError    : in     vl_logic_vector(0 to 1);
        ICU_isBus       : in     vl_logic_vector(0 to 63);
        ICU_isCA        : in     vl_logic;
        ICU_sleepReq    : in     vl_logic;
        ICU_sprDataBus  : in     vl_logic_vector(0 to 31);
        ICU_syncAfterReset: in     vl_logic;
        ICU_traceEnable : in     vl_logic;
        JTG_c405BndScanTDO: in     vl_logic;
        JTG_c405TCK     : in     vl_logic;
        JTG_c405TDI     : in     vl_logic;
        JTG_c405TMS     : in     vl_logic;
        JTG_c405TRST_NEG: in     vl_logic;
        LSSD_coreScanIn : in     vl_logic_vector(10 to 31);
        LSSD_coreTestEn : in     vl_logic;
        LSSD_jtgCClk    : in     vl_logic;
        MMU_BMCO        : in     vl_logic;
        MMU_dsStateBorC : in     vl_logic;
        MMU_dsStatus    : in     vl_logic_vector(0 to 7);
        MMU_isStatus    : in     vl_logic_vector(0 to 1);
        MMU_sprDataBus  : in     vl_logic_vector(0 to 31);
        MMU_tlbSXHit    : in     vl_logic;
        MMU_wbHold      : in     vl_logic;
        OCM_DOF         : in     vl_logic;
        OCM_dsComplete  : in     vl_logic;
        OCM_dsData      : in     vl_logic_vector(0 to 31);
        PGM_coprocPresent: in     vl_logic;
        PGM_dcu_DOF     : in     vl_logic;
        PGM_deterministicMult: in     vl_logic;
        PGM_divEn       : in     vl_logic;
        PGM_mmuEn       : in     vl_logic;
        PGM_pvrBus      : in     vl_logic_vector(0 to 31);
        PLB_dcuErr      : in     vl_logic;
        RST_c405ResetChip: in     vl_logic;
        RST_c405ResetSystem: in     vl_logic;
        TRC_c405TE      : in     vl_logic;
        TRC_c405TraceDisable: in     vl_logic;
        XXX_dcrAck      : in     vl_logic;
        XXX_dcrDataBus  : in     vl_logic_vector(0 to 31);
        XXX_uncondEvent : in     vl_logic;
        c2Clk           : in     vl_logic;
        resetCore       : in     vl_logic;
        EXE_gprSysClkPI : in     vl_logic
    );
end p405s_cpu_top;
