library verilog;
use verilog.vl_types.all;
entity p405s_DCU_logic is
    port(
        SDQ_E1          : out    vl_logic;
        SDQ_E2          : out    vl_logic;
        DCU_CA          : out    vl_logic;
        tagIndex_E1     : out    vl_logic;
        twoFP_In        : out    vl_logic;
        CAR_mmuAttr_E1  : out    vl_logic;
        CAR_mmuAttr_E2  : out    vl_logic;
        dataIndexMuxSel : out    vl_logic_vector(0 to 1);
        forceDataIndexZero_mmu: out    vl_logic;
        dataIndexMuxSel2: out    vl_logic;
        dataIndex_E2    : out    vl_logic;
        xltValidLth_E2  : out    vl_logic;
        LRU_sel0        : out    vl_logic;
        newValidIn      : out    vl_logic;
        FAR_E2          : out    vl_logic;
        newDirtyIn      : out    vl_logic;
        DCU_U0Attr_In   : out    vl_logic;
        tagIndexDup_E1  : out    vl_logic;
        tagIndexDup_E2  : out    vl_logic;
        writeTagA0      : out    vl_logic;
        dirtyLRU_readIndexSel: out    vl_logic;
        writeDataA0     : out    vl_logic;
        writeDataA1     : out    vl_logic;
        writeDirtyA0    : out    vl_logic;
        writeDirtyB0    : out    vl_logic;
        dOutMuxSelBit1Byte0: out    vl_logic;
        LRU_sel1        : out    vl_logic;
        dOutMuxSelBit1Byte1: out    vl_logic;
        dOutMuxSelBit1Byte2: out    vl_logic;
        dOutMuxSelBit1Byte3: out    vl_logic;
        flush2ndRead_In : out    vl_logic;
        FDR_lo_E2       : out    vl_logic;
        storeWord_In    : out    vl_logic;
        carFullIn       : out    vl_logic;
        storeWriting_In : out    vl_logic;
        past1stCycXltValid_In: out    vl_logic;
        writeBufMuxSelBit0: out    vl_logic;
        WB_lineDirtyIn  : out    vl_logic;
        wrAckCnt_In0X   : out    vl_logic_vector(0 to 2);
        writeBufHi_E2   : out    vl_logic_vector(0 to 3);
        CAR_OF_E2       : out    vl_logic;
        writeDirtyB1    : out    vl_logic;
        CAR_OF_full_In0 : out    vl_logic;
        FDR_hi_E1       : out    vl_logic;
        FDR_hi_E2       : out    vl_logic;
        FDR_lo_E1       : out    vl_logic;
        cacheOpMuxSel   : out    vl_logic;
        resetIn         : out    vl_logic;
        FDR_hiMuxSel    : out    vl_logic;
        FDR_holdMuxSel  : out    vl_logic;
        flushHold_E2    : out    vl_logic;
        SDP_FDR_muxSel  : out    vl_logic;
        wrAckQ_full_Inx1: out    vl_logic;
        PLBDR_hiMuxSel  : out    vl_logic_vector(0 to 3);
        wrAckQ_full_In10: out    vl_logic;
        wrAckQ_sizeTran_E1: out    vl_logic;
        wrAckQ_full_In00: out    vl_logic;
        bypassMuxSel    : out    vl_logic_vector(0 to 2);
        fillBufMuxSel0  : out    vl_logic_vector(0 to 31);
        sel_CAR_OF_full : out    vl_logic;
        fillValid_In    : out    vl_logic_vector(0 to 31);
        LSA_E2          : out    vl_logic;
        fillSM_In       : out    vl_logic_vector(0 to 5);
        FAR_full_In     : out    vl_logic;
        FAR_loadPending_In: out    vl_logic;
        dVQ_In11        : out    vl_logic_vector(0 to 6);
        PLBAR_selSAQ    : out    vl_logic;
        PLBAR_E2        : out    vl_logic;
        writeDirtyA1    : out    vl_logic;
        oneFP_In        : out    vl_logic;
        fillBuf_E2      : out    vl_logic_vector(0 to 7);
        LSA_SM_In       : out    vl_logic;
        CAR_OF_PLB_loaded_In: out    vl_logic;
        DCU_request_In  : out    vl_logic;
        xltValidLth     : out    vl_logic;
        SAQvalidNeedingPLB0: out    vl_logic;
        storeHitPend_In0: out    vl_logic_vector(0 to 1);
        SAQ_E2          : out    vl_logic;
        dirtyLRU_writeIndex_E1: out    vl_logic;
        writeTagB0      : out    vl_logic;
        DCU_sleepReq    : out    vl_logic;
        byteWriteData   : out    vl_logic_vector(0 to 15);
        dValidCnt1_In   : out    vl_logic_vector(0 to 2);
        wrAckCnt1_In    : out    vl_logic_vector(0 to 2);
        dValidCntDone_In: out    vl_logic;
        wrAckCntDone_In : out    vl_logic;
        fillFlushToDo_In: out    vl_logic;
        twoLoadPending_0_In: out    vl_logic;
        fillLineDirty_In: out    vl_logic;
        tagIndexSel     : out    vl_logic;
        dcbzFillHit_In  : out    vl_logic;
        PLBAR_E1        : out    vl_logic;
        SDQ_SDP_mux     : out    vl_logic;
        LSA_load_In     : out    vl_logic;
        priority_In     : out    vl_logic;
        DCU_guarded_In  : out    vl_logic;
        DCU_RNW_In      : out    vl_logic;
        dcbzFillHitA_In : out    vl_logic;
        writeBufLoTag_E1: out    vl_logic;
        DCU_tranSize_In : out    vl_logic;
        DCU_cacheable_In: out    vl_logic;
        SAQ_E1          : out    vl_logic;
        DCU_plbAddrBus_In: out    vl_logic_vector(30 to 31);
        cacheOpByteEn_E2: out    vl_logic;
        DCU_writeThru_In: out    vl_logic;
        cmdInProg_E2    : out    vl_logic;
        dirtyLRU_readIndex_E1: out    vl_logic;
        SAQvalidNeedingPLB1: out    vl_logic;
        DCU_byteEn_In   : out    vl_logic_vector(0 to 7);
        ocmAbort        : out    vl_logic;
        ocmLoadReq      : out    vl_logic;
        ocmStoreReq     : out    vl_logic;
        bypassFillSDP_sel: out    vl_logic_vector(0 to 3);
        dcu_DA_sel      : out    vl_logic;
        DCU_ocmWait_In0 : out    vl_logic;
        carSpecialOp_In : out    vl_logic;
        writeBufHi_E1   : out    vl_logic;
        caEarly_0_In    : out    vl_logic;
        DCUbypassPending_In0: out    vl_logic;
        cacheableSpecialOp: out    vl_logic;
        DCU_someBusy_In : out    vl_logic;
        fill_A_In       : out    vl_logic;
        carTwoFP_In     : out    vl_logic;
        LSA_bypassPending_In: out    vl_logic;
        cacheOpByteEn_E1: out    vl_logic;
        FDR_outMuxSel   : out    vl_logic_vector(0 to 1);
        carRead_In      : out    vl_logic;
        fillUsingArray  : out    vl_logic;
        CAR_OF_E1       : out    vl_logic;
        fillBufMuxSel1  : out    vl_logic_vector(0 to 31);
        PLBAR_selFAR    : out    vl_logic;
        writeBufMuxSelBit1: out    vl_logic_vector(0 to 31);
        tagOutMuxSelFAR : out    vl_logic;
        specialOPDone_In: out    vl_logic;
        fillBuf_E1      : out    vl_logic;
        specialCase_In  : out    vl_logic;
        tagReadWriteCycle_In: out    vl_logic;
        writeLRU1       : out    vl_logic;
        tagReadNotWrite_In: out    vl_logic;
        dataReadWriteCycle_In: out    vl_logic;
        carDcbzCmd      : out    vl_logic;
        DCU_firstCycCarStXltV: out    vl_logic;
        PLBDR_E2        : out    vl_logic_vector(0 to 3);
        writeTagB1      : out    vl_logic;
        dVQ_In00        : out    vl_logic_vector(0 to 6);
        dVQ_In01        : out    vl_logic_vector(0 to 6);
        LSA_E1          : out    vl_logic;
        dVQ_In10        : out    vl_logic_vector(0 to 6);
        FDR_loMuxSel    : out    vl_logic;
        LRU_out_NEG     : out    vl_logic;
        writeLRU0       : out    vl_logic;
        writeDataB0     : out    vl_logic;
        writeDataB1     : out    vl_logic;
        dataReadNotWrite_In: out    vl_logic;
        writeTagA1      : out    vl_logic;
        DCU_ocmWait_In1 : out    vl_logic;
        dcu_DA_early_NEG: out    vl_logic;
        readLRUDirty    : out    vl_logic;
        wrAckSelInc2_11 : out    vl_logic;
        setDValidCntIdle: out    vl_logic;
        wrAckCnt2_In    : out    vl_logic_vector(0 to 2);
        dValidCnt2_In   : out    vl_logic_vector(0 to 2);
        dValidCntSel    : out    vl_logic_vector(0 to 1);
        wrAckSelInc2_10 : out    vl_logic;
        DCUbypassPending_In1: out    vl_logic;
        set_storeHitPend1: out    vl_logic_vector(0 to 1);
        byteWrite_E1    : out    vl_logic;
        dataIndex_E1    : out    vl_logic;
        dirtyLRU_readIndex_E2: out    vl_logic;
        DCU_pclOcmLdPendNoWait: out    vl_logic;
        SDQ_SDP_OCM_sel : out    vl_logic;
        writeBufLo_E2   : out    vl_logic;
        storeHitFillBufPend_In: out    vl_logic;
        dataIndexLSA_dupSel: out    vl_logic;
        loadReadFBvalid : out    vl_logic;
        bypassPendOrDcRead: out    vl_logic;
        twoLoadPending_1_In: out    vl_logic;
        caEarly_1_In    : out    vl_logic;
        fillFollowedByFill_In: out    vl_logic;
        carDcRead       : out    vl_logic;
        flushIdle_state : out    vl_logic;
        flushAlmostDone : out    vl_logic;
        flushDone       : out    vl_logic;
        ocmCompleteXltVNoWaitNoHold: out    vl_logic;
        CAR_OF_fullL2   : in     vl_logic;
        dcbzFillHitA_L2 : in     vl_logic;
        fillFlushToDoL2 : in     vl_logic;
        past1stCycXltValidL2: in     vl_logic;
        carFullL2       : in     vl_logic;
        dVQ0_sizeL2     : in     vl_logic;
        fillSM          : in     vl_logic_vector(0 to 5);
        storeWritingL2  : in     vl_logic;
        xltValidL2      : in     vl_logic;
        VCT_exeAbort    : in     vl_logic;
        VCT_wbAbort     : in     vl_logic;
        storeHitPendDupL2: in     vl_logic_vector(0 to 1);
        MMU_dcuShadowAbort: in     vl_logic;
        CAR_cacheableBuf1: in     vl_logic;
        fill_A_L2       : in     vl_logic;
        SAQ_byteEn      : in     vl_logic_vector(0 to 3);
        storeHitPendL2  : in     vl_logic_vector(0 to 1);
        carOF_U0AttrL2  : in     vl_logic;
        dcbzFillHitL2   : in     vl_logic;
        ICU_dcuCCR0_L2  : in     vl_logic_vector(0 to 10);
        twoLoadPendingL2L2: in     vl_logic;
        carOF_LSAcmp    : in     vl_logic;
        U0AttrFAR       : in     vl_logic;
        carOF_FARcmp    : in     vl_logic;
        PCL_dcuOp       : in     vl_logic_vector(0 to 11);
        cacheOpBusL2    : in     vl_logic_vector(0 to 9);
        carOF_loadL2    : in     vl_logic;
        carOF_storeL2   : in     vl_logic;
        carOF_dcbzCmdL2 : in     vl_logic;
        carOF_dcbtL2    : in     vl_logic;
        carOF_cacheableL2: in     vl_logic;
        carOF_writeThruL2: in     vl_logic;
        carOF_hitAL2    : in     vl_logic;
        carOF_hitBL2    : in     vl_logic;
        carOF_byteEn    : in     vl_logic_vector(0 to 3);
        OCM_dsComplete  : in     vl_logic;
        resetL2         : in     vl_logic;
        validA          : in     vl_logic;
        validB          : in     vl_logic;
        LRU             : in     vl_logic;
        specialCaseL2   : in     vl_logic;
        dirtyA          : in     vl_logic;
        dirtyB          : in     vl_logic;
        hit_a           : in     vl_logic;
        hit_b           : in     vl_logic;
        WB_lineDirtyReadL2: in     vl_logic;
        fillLineDirtyL2 : in     vl_logic;
        CAR_writethru   : in     vl_logic;
        SAQ_L2          : in     vl_logic_vector(27 to 29);
        CAR_L2_buf1     : in     vl_logic_vector(27 to 29);
        dValidCntDoneL2 : in     vl_logic;
        wrAckCntDoneL2  : in     vl_logic;
        wrAckCntL2      : in     vl_logic_vector(0 to 2);
        carOF_dsHoldL2  : in     vl_logic;
        PLB_dcuSsizeBuf1: in     vl_logic;
        PLB_dcuWrDAck   : in     vl_logic;
        LSA_cacheableL2 : in     vl_logic;
        DCU_tranSize    : in     vl_logic;
        storeWordL2     : in     vl_logic;
        resetSCL2       : in     vl_logic;
        DCU_plbRNW_dupL2: in     vl_logic;
        LSA_L2          : in     vl_logic_vector(27 to 29);
        dVQ1_fullL2     : in     vl_logic;
        CAR_OF_L2       : in     vl_logic_vector(27 to 29);
        fillValidL2     : in     vl_logic_vector(0 to 31);
        PLB_dcuRdDAck   : in     vl_logic;
        FAR_fullL2      : in     vl_logic;
        FAR_loadPendingL2: in     vl_logic;
        PLB_dcuRdWdAddr : in     vl_logic_vector(0 to 2);
        oneFPL2         : in     vl_logic;
        LSA_SM          : in     vl_logic;
        CAR_OF_PLB_loadedL2: in     vl_logic;
        DCU_requestDupL2: in     vl_logic;
        SAQ_writeThruL2 : in     vl_logic;
        dVQ1_lineL2     : in     vl_logic;
        SAQvalidNeedingPLBL2: in     vl_logic;
        dValidCntL2     : in     vl_logic_vector(0 to 2);
        twoLoadPendingL2: in     vl_logic;
        sampleCycleL2   : in     vl_logic;
        carByteEn       : in     vl_logic_vector(0 to 3);
        twoFPL2         : in     vl_logic;
        LSA_loadL2      : in     vl_logic;
        CAR_LSAcmp      : in     vl_logic;
        dVQ1_sizeL2     : in     vl_logic;
        SAQ_cacheableL2 : in     vl_logic;
        ICU_syncAfterReset: in     vl_logic;
        dVQ0_fullL2     : in     vl_logic_vector(0 to 1);
        carOF_guardedL2 : in     vl_logic;
        SAQ_FARcmp      : in     vl_logic;
        wrAckQ_sizeL2   : in     vl_logic;
        SAQ_guardedL2   : in     vl_logic;
        SAQ_U0AttrL2    : in     vl_logic;
        DCU_someBusyL2  : in     vl_logic;
        OCM_dsHold      : in     vl_logic;
        MMU_wbHold      : in     vl_logic;
        CAR_SAQcmp      : in     vl_logic;
        carSpecialOpL2  : in     vl_logic;
        caEarlyL2       : in     vl_logic;
        DCUbypassPendingL2: in     vl_logic;
        DCU_ocmWait     : in     vl_logic;
        dVQ0_lineL2     : in     vl_logic;
        busySCL2        : in     vl_logic;
        wrAckQ_fullL2   : in     vl_logic;
        wrAckQ_lineL2   : in     vl_logic;
        carTwoFPL2      : in     vl_logic;
        LSA_bypassPendingL2: in     vl_logic;
        carReadL2       : in     vl_logic;
        resetCore       : in     vl_logic;
        specialOPDoneL2 : in     vl_logic;
        MMU_dcuUTLBAbortL2: in     vl_logic;
        flush2ndReadL2  : in     vl_logic;
        storeHitFillBufPendL2: in     vl_logic;
        PLB_dcuRdDAck2  : in     vl_logic;
        dValidCntDone2L2: in     vl_logic;
        fillSM2         : in     vl_logic_vector(0 to 5);
        CAR_OF_full2L2  : in     vl_logic;
        CAR_cacheableBuf2: in     vl_logic;
        reset4L2        : in     vl_logic;
        PCL_dcuOp_early : in     vl_logic_vector(0 to 2);
        CAR_cacheableNoBuf: in     vl_logic;
        xltValidDupL2   : in     vl_logic;
        testEn          : in     vl_logic;
        LSA_guardedL2   : in     vl_logic;
        carFull2L2      : in     vl_logic;
        fillFollowedByFillL2: in     vl_logic;
        PLB_dcuWrDAckBuf: in     vl_logic;
        PLB_dcuRdDAck3  : in     vl_logic;
        carLoadDup      : in     vl_logic;
        carStoreDup     : in     vl_logic;
        CAR_L2_buf2     : in     vl_logic_vector(27 to 29);
        PLB_dcuSsizeBuf2: in     vl_logic;
        SAQvalidNeedingPLB2L2: in     vl_logic;
        fillSM3_pend    : in     vl_logic;
        dValidCntDone3L2: in     vl_logic
    );
end p405s_DCU_logic;
