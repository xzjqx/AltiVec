library verilog;
use verilog.vl_types.all;
entity p405s_icu_ram_data_flow_16K is
    port(
        ICU_isBus       : out    vl_logic_vector(0 to 63);
        ICU_parityErrE  : out    vl_logic;
        ICU_parityErrO  : out    vl_logic;
        ICU_tagParityErr: out    vl_logic;
        compareA        : out    vl_logic;
        compareA_NEG    : out    vl_logic;
        compareB        : out    vl_logic;
        compareB_NEG    : out    vl_logic;
        dsCompA         : out    vl_logic;
        dsCompB         : out    vl_logic;
        icReadData      : out    vl_logic_vector(0 to 31);
        icuCacheSize    : out    vl_logic_vector(0 to 2);
        lruOut          : out    vl_logic;
        vaOut           : out    vl_logic;
        vbOut           : out    vl_logic;
        CB              : in     vl_logic;
        ICU_paritySel   : in     vl_logic;
        ICU_baSel       : in     vl_logic;
        ICU_tagDataSel  : in     vl_logic;
        JTG_iCacheWr    : in     vl_logic;
        JTG_inst        : in     vl_logic_vector(0 to 31);
        Lx27Sel         : in     vl_logic;
        Lx28Sel         : in     vl_logic;
        Lx29Sel         : in     vl_logic;
        MMU_isCacheable : in     vl_logic;
        MMU_isRA        : in     vl_logic_vector(0 to 21);
        OCM_isData      : in     vl_logic_vector(0 to 63);
        PLB_icuDBus     : in     vl_logic_vector(0 to 63);
        VaVbRdSel       : in     vl_logic_vector(0 to 2);
        VaVbWrE1        : in     vl_logic;
        cycleDataRegAIn : in     vl_logic;
        cycleDataRegBIn : in     vl_logic;
        cycleTagRegIn   : in     vl_logic;
        cycleParityRegIn: in     vl_logic;
        dataRdWrRegIn   : in     vl_logic;
        df_dataCc       : in     vl_logic_vector(18 to 27);
        df_jtagIsEa_NEG : in     vl_logic_vector(18 to 26);
        df_lruRdCcInNEG : in     vl_logic_vector(18 to 26);
        df_lruWrCcIn    : in     vl_logic_vector(18 to 26);
        df_rars         : in     vl_logic_vector(0 to 21);
        df_rarsTLE      : in     vl_logic;
        df_tagVccRegIn  : in     vl_logic_vector(18 to 26);
        dsRD1cycle      : in     vl_logic;
        fillAE2         : in     vl_logic_vector(0 to 7);
        fillBE2         : in     vl_logic_vector(0 to 7);
        fillWr0L2       : in     vl_logic;
        isBusSel        : in     vl_logic_vector(0 to 1);
        lruRdCcE1       : in     vl_logic;
        newLruBitIn     : in     vl_logic;
        newVaBitIn      : in     vl_logic;
        newVbBitIn      : in     vl_logic;
        rdStateL2       : in     vl_logic;
        rdar            : in     vl_logic_vector(0 to 29);
        scL2            : in     vl_logic;
        tagBWE1         : in     vl_logic;
        tagRdWrRegIn    : in     vl_logic;
        vaOutL2         : in     vl_logic;
        vbOutL2         : in     vl_logic;
        wbHighE2        : in     vl_logic_vector(0 to 3);
        wbLowE2         : in     vl_logic;
        wbTagE1         : in     vl_logic;
        wrATagNotB      : in     vl_logic;
        wrFlashIn       : in     vl_logic;
        wrLruIn         : in     vl_logic_vector(0 to 2);
        wrVaIn          : in     vl_logic;
        wrVbIn          : in     vl_logic;
        ICU_CCR1ICTE    : in     vl_logic;
        ICU_CCR1ICDE    : in     vl_logic;
        resetMemBist    : in     vl_logic;
        icu_bist_debug_si: in     vl_logic_vector(3 downto 0);
        icu_bist_debug_so: out    vl_logic_vector(3 downto 0);
        icu_bist_debug_en: in     vl_logic_vector(3 downto 0);
        icu_bist_mode_reg_in: in     vl_logic_vector(18 downto 0);
        icu_bist_mode_reg_out: out    vl_logic_vector(18 downto 0);
        icu_bist_parallel_dr: in     vl_logic;
        icu_bist_mode_reg_si: in     vl_logic;
        icu_bist_mode_reg_so: out    vl_logic;
        icu_bist_shift_dr: in     vl_logic;
        icu_bist_mbrun  : in     vl_logic
    );
end p405s_icu_ram_data_flow_16K;
