library verilog;
use verilog.vl_types.all;
entity p405s_icu_hitPath is
    port(
        BufValidIn_NEG  : out    vl_logic;
        ICU_mmuEoOdd    : out    vl_logic;
        ICU_ocmIcuReady_NEG: out    vl_logic;
        VaVbRdSel       : out    vl_logic_vector(0 to 2);
        compAlru_NEG    : out    vl_logic;
        compB_NEG       : out    vl_logic;
        cycleDataRegAIn : out    vl_logic;
        cycleDataRegBIn : out    vl_logic;
        cycleParityRegIn: out    vl_logic;
        cycleTagRegIn   : out    vl_logic;
        eo_0            : out    vl_logic;
        eo_1            : out    vl_logic;
        forceNlIn       : out    vl_logic;
        lxFetchValidIn  : out    vl_logic;
        lxSel           : out    vl_logic;
        missIn          : out    vl_logic;
        nxtFetchRd      : out    vl_logic;
        nxtWait         : out    vl_logic;
        rdStateIn       : out    vl_logic;
        tagVSel_0       : out    vl_logic;
        vcarSelHi_NEG   : out    vl_logic;
        vcarSelLow_NEG  : out    vl_logic;
        vcarSel_pri_NEG : out    vl_logic;
        wrLruIn         : out    vl_logic_vector(0 to 2);
        IFB_isAbort2    : in     vl_logic;
        IFB_isNL        : in     vl_logic;
        OCM_isHold      : in     vl_logic;
        VaVb_VR_pg4_NEG : in     vl_logic;
        bufValidL2_NEG  : in     vl_logic;
        compareA        : in     vl_logic;
        compareA_NEG    : in     vl_logic;
        compareB        : in     vl_logic;
        compareB_NEG    : in     vl_logic;
        cycle_RA_p3_NEG : in     vl_logic;
        cycle_RB_p3_NEG : in     vl_logic;
        cycle_parity_p3_NEG: in     vl_logic;
        cycle_RT_p3_NEG : in     vl_logic;
        eo_q            : in     vl_logic;
        eo_r            : in     vl_logic;
        eo_y_NEG        : in     vl_logic;
        eo_z2_NEG       : in     vl_logic;
        eo_z_NEG        : in     vl_logic;
        forceNlL2       : in     vl_logic;
        frAndDsRdy      : in     vl_logic;
        ldcc2RdNoAb_NEG : in     vl_logic;
        lxFetchValidIn_A_NEG: in     vl_logic;
        lxFetchValidIn_B_NEG: in     vl_logic;
        lxFetchValidL2  : in     vl_logic;
        lxSel_C_NEG     : in     vl_logic;
        lxSel_D_NEG     : in     vl_logic;
        missL2          : in     vl_logic;
        nfr_ABC_p2_NEG  : in     vl_logic;
        nxtWa_W_NEG     : in     vl_logic;
        nxtWa_X_NEG     : in     vl_logic;
        ocmDvQ_1_NEG    : in     vl_logic;
        rdOrWaAndXltValid: in     vl_logic;
        rdSt_RDA_pg4_NEG: in     vl_logic;
        setForceNl      : in     vl_logic;
        tagSelBit0_E_NEG: in     vl_logic;
        tagSelBit0_F_NEG: in     vl_logic;
        vcarSel_noEO    : in     vl_logic;
        wrLruNoHit_NEG  : in     vl_logic
    );
end p405s_icu_hitPath;
