library verilog;
use verilog.vl_types.all;
entity p405s_exeStage is
    port(
        PCL_dcuOp       : out    vl_logic_vector(0 to 11);
        PCL_dsMmuOp     : out    vl_logic_vector(0 to 3);
        PCL_exeAdmCntl  : out    vl_logic_vector(0 to 3);
        PCL_exeCmplmntA : out    vl_logic;
        PCL_exeApuOp    : out    vl_logic;
        PCL_exeCpuOp    : out    vl_logic;
        PCL_exeWrExtEn  : out    vl_logic;
        PCL_exeLogicalCntl: out    vl_logic_vector(0 to 7);
        PCL_exePrivOp   : out    vl_logic;
        PCL_exeSprDataEn_NEG: out    vl_logic;
        PCL_exeSrmCntl  : out    vl_logic_vector(0 to 3);
        PCL_exeXerCaEn  : out    vl_logic;
        PCL_exeXerOvEn  : out    vl_logic;
        PCL_icuOp       : out    vl_logic_vector(0 to 3);
        PCL_ldNotSt     : out    vl_logic;
        PCL_mfSPR       : out    vl_logic;
        PCL_mtSPR       : out    vl_logic;
        PCL_nopStringIndexed: out    vl_logic;
        PCL_tlbRE       : out    vl_logic;
        PCL_tlbSX       : out    vl_logic;
        PCL_tlbWE       : out    vl_logic;
        PCL_tlbWS       : out    vl_logic;
        exeFull         : out    vl_logic;
        exeLSSMIURA     : out    vl_logic_vector(0 to 7);
        exeMfdcr        : out    vl_logic;
        exeMtdcr        : out    vl_logic;
        exeRpWrEn       : out    vl_logic;
        exeXerTBCUpdInstr: out    vl_logic;
        APU_dcdPrivOp   : in     vl_logic;
        CB              : in     vl_logic;
        EXE_xerTBCNotEqZero: in     vl_logic;
        APU_dcdApuOp    : in     vl_logic;
        plaVal          : in     vl_logic;
        dcdRegBit20     : in     vl_logic;
        dcdXerTBCUpdInstr: in     vl_logic;
        exeClearOrFlush : in     vl_logic;
        exeE1           : in     vl_logic;
        exeE2           : in     vl_logic;
        gtErr           : in     vl_logic;
        plaAdmCntl      : in     vl_logic_vector(0 to 3);
        plaAddEn        : in     vl_logic;
        plaCmplmntA     : in     vl_logic;
        plaDcuOp        : in     vl_logic_vector(0 to 11);
        plaEaCalc       : in     vl_logic;
        plaIcuOp        : in     vl_logic_vector(0 to 3);
        plaWrExtEn      : in     vl_logic;
        plaLSSMIURA     : in     vl_logic_vector(0 to 7);
        plaLdNotSt      : in     vl_logic;
        plaLogicalCntl  : in     vl_logic_vector(0 to 7);
        plaMfdcr        : in     vl_logic;
        plaMfspr        : in     vl_logic;
        plaMmuCode      : in     vl_logic_vector(0 to 6);
        plaMtdcr        : in     vl_logic;
        plaMtspr        : in     vl_logic;
        plaOeCk         : in     vl_logic;
        plaPriv         : in     vl_logic;
        plaRpWrEn       : in     vl_logic;
        plaSrmCntl      : in     vl_logic_vector(0 to 3);
        plaUnitEn       : in     vl_logic_vector(0 to 4);
        plaXerCaEn      : in     vl_logic;
        nxtExeFull      : in     vl_logic;
        exeStorageOp    : out    vl_logic;
        plaLwarx        : in     vl_logic;
        plaStwcx        : in     vl_logic;
        exeLwarx        : out    vl_logic;
        exeStwcx        : out    vl_logic;
        NplaApRdEn      : in     vl_logic;
        NplaBpRdEn      : in     vl_logic;
        plaSpRdEn       : in     vl_logic;
        exeApRdEn       : out    vl_logic;
        exeBpRdEn       : out    vl_logic;
        exeSpRdEn       : out    vl_logic;
        plaWrtee        : in     vl_logic;
        PCL_exeWrtee    : out    vl_logic;
        APU_dcdLoad     : in     vl_logic;
        APU_dcdStore    : in     vl_logic;
        APU_dcdUpdate   : in     vl_logic;
        APU_dcdFpuOp    : in     vl_logic;
        exeApuFpuOp     : out    vl_logic;
        exeApuFpuLoad   : out    vl_logic;
        PCL_exe2DataE1  : in     vl_logic;
        PCL_exe2DataE2  : in     vl_logic;
        exe2ClearOrFlush: in     vl_logic;
        exe2Full        : out    vl_logic;
        PCL_exeNegMac   : out    vl_logic;
        PCL_exeFpuOp    : out    vl_logic;
        dcdApuValidOp_NEG: in     vl_logic;
        APU_dcdGprWr    : in     vl_logic;
        PCL_exeApuValidOp: out    vl_logic;
        plaMac          : in     vl_logic;
        plaNegMac       : in     vl_logic;
        exeRpEqexe2RpAddr: in     vl_logic;
        PCL_exe2AccRegMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exe2NegMac  : out    vl_logic;
        PCL_exe2MacEn   : out    vl_logic;
        PCL_exe2MultEn  : out    vl_logic;
        PCL_exe2MultHiWd: out    vl_logic;
        PCL_exe2XerOvEn : out    vl_logic;
        PCL_exeRbEn     : out    vl_logic_vector(0 to 3);
        PCL_exeDbgRdOp  : out    vl_logic;
        PCL_exeDbgWrOp  : out    vl_logic;
        APU_dcdXerCAEn  : in     vl_logic;
        APU_dcdXerOVEn  : in     vl_logic;
        dcdMmuSprDcd    : in     vl_logic_vector(0 to 8);
        PCL_mmuSprDcd   : out    vl_logic_vector(0 to 8);
        exeStrgSt       : in     vl_logic_vector(1 to 2);
        PCL_exeMultEn   : out    vl_logic;
        PCL_exeDivEn    : out    vl_logic;
        PCL_exeLogicalUnitEn_NEG: out    vl_logic;
        PCL_exeSrmUnitEn_NEG: out    vl_logic;
        PCL_exeSprUnitEn_NEG: out    vl_logic;
        exeEaCalc       : out    vl_logic;
        PCL_exeAddEn    : out    vl_logic;
        PCL_exeMacEn    : out    vl_logic;
        PCL_exeRaEn     : out    vl_logic_vector(0 to 3);
        PCL_exeStringMultiple: out    vl_logic;
        plaGateZeroToAccReg: in     vl_logic;
        dcdSecOpBit21L2 : in     vl_logic;
        dcdRSRTL2       : in     vl_logic_vector(0 to 4);
        PCL_exeTrapCond : out    vl_logic_vector(0 to 4);
        exeLoadQ        : out    vl_logic;
        plaMacSat       : in     vl_logic;
        PCL_exe2MacSat  : out    vl_logic;
        exeMmuOp        : out    vl_logic;
        PCL_Rbit        : in     vl_logic;
        plaSrmBpSel     : in     vl_logic_vector(0 to 2);
        PCL_exeSrmBpSel : out    vl_logic_vector(0 to 2);
        PCL_exe2SignedOp: out    vl_logic;
        exeMultEn       : out    vl_logic;
        exeMacEn        : out    vl_logic;
        PCL_exeDbgLdOp  : out    vl_logic;
        PCL_exeDbgStOp  : out    vl_logic;
        APU_dcdRaEn     : in     vl_logic;
        APU_dcdRbEn     : in     vl_logic;
        APU_dcdForceAlgn: in     vl_logic;
        APU_dcdExeLdDepend: in     vl_logic;
        exeDivEn        : out    vl_logic;
        APU_dcdWbLdDepend: in     vl_logic;
        APU_dcdLwbLdDepend: in     vl_logic;
        exeApuExeWbLdUseL2: out    vl_logic;
        exeApuExeLwbLdUseL2: out    vl_logic;
        PCL_exeMultEn_NEG: out    vl_logic_vector(0 to 1);
        PCL_exeDivEnForMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exeCmplmntA_NEG: out    vl_logic;
        PCL_exe2MacOrMultEn_NEG: out    vl_logic_vector(0 to 1);
        PCL_exe2MacOrMultEnForMS: out    vl_logic_vector(0 to 1);
        PCL_exeMultEnForMuxSel: out    vl_logic_vector(0 to 1);
        wbHold          : in     vl_logic;
        ltchDA          : in     vl_logic;
        PCL_exeEaCalc   : out    vl_logic;
        plaApuLdSt      : in     vl_logic;
        exeForceAlgn    : out    vl_logic;
        dcdIcuSprDcd    : in     vl_logic_vector(0 to 2);
        dcdTimSprDcd    : in     vl_logic_vector(0 to 5);
        PCL_icuSprDcds  : out    vl_logic_vector(0 to 2);
        PCL_timSprDcds  : out    vl_logic_vector(0 to 5);
        dcdDbgSprDcd    : in     vl_logic_vector(0 to 3);
        dcdExeSprDcd    : in     vl_logic_vector(0 to 4);
        dcdVctSprDcd    : in     vl_logic_vector(0 to 5);
        PCL_dbgSprDcds  : out    vl_logic_vector(0 to 3);
        PCL_exeSprDcds  : out    vl_logic_vector(0 to 4);
        PCL_vctSprDcds  : out    vl_logic_vector(0 to 5);
        resetL2         : in     vl_logic;
        plaForceAlgn    : in     vl_logic;
        PCL_exeAddSgndOp_NEG: out    vl_logic_vector(0 to 1);
        PCL_exeDivSgndOp: out    vl_logic;
        PCL_exeDivEn_NEG: out    vl_logic;
        PCL_dcuOp_early : out    vl_logic_vector(0 to 2);
        exeFullForE1_NEG: out    vl_logic;
        exe2FullForE1_NEG: out    vl_logic;
        APU_dcdTrapLE   : in     vl_logic;
        APU_dcdTrapBE   : in     vl_logic;
        APU_dcdForceBESteering: in     vl_logic;
        exeTrapLE       : out    vl_logic;
        exeTrapBE       : out    vl_logic;
        exeForceBESteering: out    vl_logic;
        PCL_exeMacOrMultEn_NEG: out    vl_logic;
        plaMtcrf        : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        PCL_exeDivEnForLSSD: out    vl_logic;
        IFB_dcdFull     : in     vl_logic;
        countE1         : out    vl_logic;
        PCL_exeSrmUnitEnForLSSD: out    vl_logic;
        exeApuFpuLdSt   : out    vl_logic;
        PCL_exeLogicalUnitEnForLSSD: out    vl_logic;
        exeStrgStC0     : in     vl_logic;
        PCL_exeTlbOp    : out    vl_logic;
        dcdJtgSprDcd    : in     vl_logic;
        PCL_jtgSprDcd   : out    vl_logic
    );
end p405s_exeStage;
