library verilog;
use verilog.vl_types.all;
entity p405s_fetcher is
    port(
        IFB_dcdApu      : out    vl_logic_vector(0 to 31);
        IFB_dcdDataIn_Neg: out    vl_logic_vector(0 to 31);
        IFB_exeDisableDbL2: out    vl_logic;
        IFB_exeIfetchErrL2: out    vl_logic_vector(0 to 4);
        IFB_iac1BitsEq  : out    vl_logic;
        IFB_iac1GtIar   : out    vl_logic;
        IFB_iac2BitsEq  : out    vl_logic;
        IFB_iac2GtIar   : out    vl_logic;
        IFB_iac3BitsEq  : out    vl_logic;
        IFB_iac3GtIar   : out    vl_logic;
        IFB_iac4BitsEq  : out    vl_logic;
        IFB_iac4GtIar   : out    vl_logic;
        IFB_isEA        : out    vl_logic_vector(0 to 29);
        IFB_isNL        : out    vl_logic;
        IFB_isNP        : out    vl_logic;
        IFB_isOcmAbus   : out    vl_logic_vector(0 to 29);
        IFB_traceData   : out    vl_logic_vector(0 to 29);
        IFB_wbDisableDbL2: out    vl_logic;
        IFB_wbIar       : out    vl_logic_vector(0 to 29);
        dcdData2L2      : out    vl_logic_vector(11 to 15);
        dcdDataBD_0     : out    vl_logic;
        dcdDataBO       : out    vl_logic_vector(0 to 4);
        dcdDataL2       : out    vl_logic_vector(0 to 31);
        dcdDataPri      : out    vl_logic_vector(0 to 5);
        dcdDataSec      : out    vl_logic_vector(0 to 10);
        exeIarL2        : out    vl_logic_vector(0 to 29);
        isEaBuf         : out    vl_logic_vector(0 to 29);
        lcar_29         : out    vl_logic;
        pfb0DataL2      : out    vl_logic_vector(0 to 31);
        refetchPipeAddr : out    vl_logic_vector(0 to 29);
        wbBrTakenL2     : out    vl_logic;
        wbTEL2          : out    vl_logic_vector(0 to 4);
        CB              : in     vl_logic;
        DBG_exeTE       : in     vl_logic_vector(0 to 4);
        DBG_iacEn       : in     vl_logic;
        ICU_ifbEDataBus : in     vl_logic_vector(0 to 31);
        ICU_ifbError    : in     vl_logic_vector(0 to 1);
        ICU_ifbODataBus : in     vl_logic_vector(0 to 31);
        IFB_exeDbgBrTaken: in     vl_logic;
        JTG_dbdrPulse   : in     vl_logic;
        JTG_inst        : in     vl_logic_vector(0 to 31);
        LSSD_coreTestEn : in     vl_logic;
        MMU_isStatus    : in     vl_logic_vector(0 to 1);
        PCL_exe2Full    : in     vl_logic;
        PCL_exe2IarE1   : in     vl_logic;
        PCL_exe2IarE2   : in     vl_logic;
        VCT_vectorBus   : in     vl_logic_vector(0 to 7);
        coreResetL2     : in     vl_logic;
        ctrL2           : in     vl_logic_vector(0 to 29);
        dbsrPulseCntlE1 : in     vl_logic;
        dcdApuE1        : in     vl_logic;
        dcdBrTarSel     : in     vl_logic_vector(0 to 1);
        dcdCorrect_Neg  : in     vl_logic;
        dcdCrtBpntLrCtr : in     vl_logic;
        dcdCrtE2        : in     vl_logic;
        dcdCrtMuxSel    : in     vl_logic;
        dcdDataMuxSel   : in     vl_logic_vector(0 to 1);
        dcdE1           : in     vl_logic;
        dcdE2           : in     vl_logic;
        dcdFullL2       : in     vl_logic;
        dcdIarMuxSel    : in     vl_logic_vector(0 to 1);
        dcdTarget_Neg   : in     vl_logic;
        evprL2          : in     vl_logic_vector(0 to 15);
        exeCorrect_Neg  : in     vl_logic;
        exeCrtBpntLrCtr : in     vl_logic;
        exeCrtE2        : in     vl_logic;
        exeCrtMuxSel    : in     vl_logic_vector(0 to 1);
        exeDataBr_21L2  : in     vl_logic;
        exeDataE1       : in     vl_logic;
        exeDataE2       : in     vl_logic;
        exeFlushorClear : in     vl_logic;
        exeIarE2        : in     vl_logic;
        iac1L2          : in     vl_logic_vector(0 to 29);
        iac2L2          : in     vl_logic_vector(0 to 29);
        iac3L2          : in     vl_logic_vector(0 to 29);
        iac4L2          : in     vl_logic_vector(0 to 29);
        isEaMuxSel      : in     vl_logic;
        isEa_22DlyL2    : in     vl_logic;
        isEa_27DlyL2    : in     vl_logic;
        lcarE2          : in     vl_logic;
        lcarMuxSel      : in     vl_logic_vector(0 to 1);
        linkL2          : in     vl_logic_vector(0 to 29);
        lrCtrNormal_Neg : in     vl_logic_vector(0 to 29);
        lrCtrSe_Neg     : in     vl_logic_vector(0 to 29);
        mux048Sel       : in     vl_logic_vector(0 to 1);
        pfb0BrTarSel    : in     vl_logic_vector(0 to 1);
        pfb0DataMuxSel  : in     vl_logic_vector(0 to 1);
        pfb0E1          : in     vl_logic;
        pfb0E2          : in     vl_logic;
        pfb0IarMuxSel   : in     vl_logic_vector(0 to 1);
        pfb1DataMuxSel  : in     vl_logic;
        pfb1E2          : in     vl_logic;
        pfb1IarMuxSel   : in     vl_logic;
        refetchAddrSel  : in     vl_logic;
        refetchLcarMuxSel: in     vl_logic_vector(0 to 1);
        refetchPipeStageSel: in     vl_logic_vector(0 to 1);
        saveForTraceE1  : in     vl_logic;
        saveForTraceE2  : in     vl_logic;
        srr02_Neg       : in     vl_logic_vector(0 to 29);
        traceDataSel    : in     vl_logic_vector(0 to 1);
        tracePipeStageSel: in     vl_logic_vector(0 to 1);
        wbDataE1        : in     vl_logic;
        wbDataE2        : in     vl_logic;
        wbFlushOrClear  : in     vl_logic;
        wbIarE1         : in     vl_logic;
        wbIarE2         : in     vl_logic;
        MMU_isParityErr : in     vl_logic;
        ICU_parityErrE  : in     vl_logic;
        ICU_tagParityErr: in     vl_logic;
        ICU_parityErrO  : in     vl_logic;
        IFB_exeISideMachChk: out    vl_logic;
        ICU_CCR0IPE     : in     vl_logic;
        ICU_CCR0TPE     : in     vl_logic
    );
end p405s_fetcher;
