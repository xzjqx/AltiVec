library verilog;
use verilog.vl_types.all;
entity p405s_admCntl is
    port(
        EXE_admMco      : out    vl_logic;
        aRegMuxSel      : out    vl_logic_vector(0 to 1);
        admOutMuxSel    : out    vl_logic_vector(0 to 1);
        multLoAnsMuxSel : out    vl_logic;
        bRegMuxSel      : out    vl_logic_vector(0 to 1);
        sgndOpNotZero   : out    vl_logic;
        dndSE_NEG       : out    vl_logic;
        sRegMuxSel      : out    vl_logic_vector(0 to 1);
        addOV           : out    vl_logic;
        divOV           : out    vl_logic;
        nxtQ            : out    vl_logic;
        PCL_aPortRregBypass: in     vl_logic;
        PCL_bPortRregBypass: in     vl_logic;
        PCL_exeCmplmntA : in     vl_logic;
        PCL_dcdHotCIn   : in     vl_logic;
        PCL_dcdXerCa    : in     vl_logic;
        PCL_exeDivEn    : in     vl_logic;
        PCL_exeMultEn   : in     vl_logic;
        PCL_sPortRregBypass: in     vl_logic;
        N_ZP            : in     vl_logic;
        aBytes01Eq0     : in     vl_logic;
        bBytes23Eq0     : in     vl_logic;
        adderOutBit0    : in     vl_logic;
        adderOutBit16   : in     vl_logic;
        adderOutSgnBit  : in     vl_logic;
        coreReset       : in     vl_logic;
        deterministicMult: in     vl_logic;
        divSt           : in     vl_logic_vector(0 to 5);
        bBusBit0        : in     vl_logic;
        sBusBit0        : in     vl_logic;
        bBytes01Eq0     : in     vl_logic;
        N_OP            : in     vl_logic;
        multHiWd        : in     vl_logic;
        nxtXerCa        : in     vl_logic;
        aBusBit0        : in     vl_logic;
        aBusBit16       : in     vl_logic;
        bBusBit16       : in     vl_logic;
        signedOp        : in     vl_logic;
        bBytes01Eq1     : in     vl_logic;
        aBytes01Eq1     : in     vl_logic;
        PCL_holdCIn     : in     vl_logic;
        PCL_gateZeroToAreg: in     vl_logic;
        PCL_gateZeroToSreg: in     vl_logic;
        PCL_addFour     : in     vl_logic;
        multSt          : in     vl_logic_vector(0 to 1);
        CB              : in     vl_logic;
        CIn             : out    vl_logic;
        PCL_dcdSrmBpSel : in     vl_logic_vector(0 to 2);
        srmMuxSel       : out    vl_logic_vector(0 to 5);
        multOV          : out    vl_logic;
        EXE_multMco     : out    vl_logic;
        divStE2         : out    vl_logic;
        multStE2        : out    vl_logic;
        PCL_wbHold      : in     vl_logic;
        multAnsLoBit0   : in     vl_logic;
        multLWAnsLoE1   : out    vl_logic;
        multLWAnsHiE1   : out    vl_logic;
        divPathEn       : out    vl_logic;
        PCL_exeXerOvEn  : in     vl_logic;
        PCL_dcdAregLoadUse: in     vl_logic;
        PCL_dcdBregLoadUse: in     vl_logic;
        PCL_dcdSregLoadUse: in     vl_logic;
        PCL_bPortLitGenSel: in     vl_logic;
        PCL_exeAregLoadUse: in     vl_logic;
        PCL_exeBregLoadUse: in     vl_logic;
        PCL_exeSregLoadUse: in     vl_logic;
        mdSgn           : out    vl_logic;
        mrSgn           : out    vl_logic;
        EXE_divMco      : out    vl_logic;
        divASeEn        : out    vl_logic;
        nonDivASeEn     : out    vl_logic;
        macMdMuxSel     : out    vl_logic;
        macMrMuxSel     : out    vl_logic;
        macRsHiEn       : out    vl_logic;
        macRsLoEn       : out    vl_logic_vector(0 to 1);
        lastCycSgnMd    : out    vl_logic;
        firstCycSgnMd   : out    vl_logic;
        exe2MacE1       : out    vl_logic;
        accRegE1        : out    vl_logic;
        PCL_dcdMrSelQ   : in     vl_logic;
        PCL_dcdMdSelQ   : in     vl_logic;
        macRcHiEn       : out    vl_logic;
        macRcLoEn       : out    vl_logic_vector(0 to 1);
        tczPSHiMuxSel   : out    vl_logic_vector(0 to 1);
        tcPSLoMuxSel    : out    vl_logic;
        tczPCHiMuxSel   : out    vl_logic_vector(0 to 1);
        tcPCLoMuxSel    : out    vl_logic;
        md2CompEn       : out    vl_logic;
        PCL_exe2MultEn  : in     vl_logic;
        PCL_exe2MultHiWd: in     vl_logic;
        PCL_exe2XerOvEn : in     vl_logic;
        PCL_exe2Hold    : in     vl_logic;
        PCL_exe2NegMac  : in     vl_logic;
        PCL_exeMacEn    : in     vl_logic;
        multCntr        : in     vl_logic_vector(0 to 1);
        nxtMultCntr     : out    vl_logic_vector(0 to 1);
        adderOutBit15   : in     vl_logic;
        divNxtToLastSt  : out    vl_logic;
        divLastStOrSt0L2: in     vl_logic;
        OPHi16          : in     vl_logic;
        ZPHi16          : in     vl_logic;
        exe2Mult16x32   : out    vl_logic;
        exe2Mult16x16Signed: out    vl_logic;
        resetL2         : out    vl_logic;
        ZPLo16          : in     vl_logic;
        OPLo16          : in     vl_logic;
        multLWAnsLo     : in     vl_logic_vector(0 to 15);
        multLWAnsHi     : in     vl_logic_vector(0 to 15);
        PCL_exeNegMac   : in     vl_logic;
        multHiEOAnsCc   : out    vl_logic_vector(0 to 2);
        multLo4CycAnsCc : out    vl_logic_vector(0 to 2);
        multLo5CycAnsCc : out    vl_logic_vector(0 to 2);
        PCL_exe2MacEn   : in     vl_logic;
        PCL_exe2MacSat  : in     vl_logic;
        macOV           : out    vl_logic;
        PCL_exeLoadUseHold: in     vl_logic;
        PCL_exeDvcHold  : in     vl_logic;
        PCL_exeSrmBpSel : in     vl_logic_vector(0 to 2);
        MDBit0          : in     vl_logic;
        MRBit0          : in     vl_logic;
        macAccL2Bit0    : in     vl_logic;
        PCL_exe2SignedOp: in     vl_logic;
        PCL_holdMdMr    : in     vl_logic;
        exe2MacE2       : out    vl_logic;
        divLastStOrSt0L2_NEG: in     vl_logic;
        macCarryBit2    : in     vl_logic;
        macSumBit1      : in     vl_logic;
        PCL_exeAddSgndOp_NEG: in     vl_logic_vector(0 to 1);
        PCL_exeDivSgndOp: in     vl_logic;
        PCL_exeDivEn_NEG: in     vl_logic;
        divSt1_NEG      : in     vl_logic;
        divSt0Or1       : in     vl_logic;
        PCL_exeDivEnForLSSD: in     vl_logic;
        cIn_1           : out    vl_logic;
        exe2MacProdSgndL2: out    vl_logic;
        exe2MacSatUnsigned: out    vl_logic;
        exe2Md16BitOprndL2: out    vl_logic;
        exe2Mr16BitOprndL2: out    vl_logic;
        potSOV          : out    vl_logic;
        sumBit1         : out    vl_logic;
        nxtQ_NEG        : out    vl_logic;
        PCL_exeDvcOrParityHold: in     vl_logic
    );
end p405s_admCntl;
