library verilog;
use verilog.vl_types.all;
entity p405s_fileAddrCntl is
    port(
        dcdRAEqlwbLpAddr: out    vl_logic;
        dcdRAEqwbLpAddr : out    vl_logic;
        dcdRAEqwbRpAddr : out    vl_logic;
        dcdRAEqexeRpAddr: out    vl_logic;
        dcdRBEqlwbLpAddr: out    vl_logic;
        dcdRBEqwbLpAddr : out    vl_logic;
        dcdRBEqwbRpAddr : out    vl_logic;
        dcdRBEqexeRpAddr: out    vl_logic;
        dcdRSEqlwbLpAddr: out    vl_logic;
        dcdRSEqwbLpAddr : out    vl_logic;
        dcdRSEqwbRpAddr : out    vl_logic;
        dcdRSEqexeRpAddr: out    vl_logic;
        dcdRAEqexeMorMRpAddr: out    vl_logic;
        dcdRBEqexeMorMRpAddr: out    vl_logic;
        dcdRSEqexeMorMRpAddr: out    vl_logic;
        exeRSEqlwbLpAddr: out    vl_logic;
        exeRSEqwbRpAddr : out    vl_logic;
        exeRpEqdcdSpAddr: out    vl_logic;
        exeRpEqwbLpAddr : out    vl_logic;
        exeRpEqlwbLpAddr: out    vl_logic;
        lwbLpEqexeApAddr: out    vl_logic;
        lwbLpEqexeBpAddr: out    vl_logic;
        lwbLpEqexeSpAddr: out    vl_logic;
        wbLpEqexeApAddr : out    vl_logic;
        wbLpEqexeBpAddr : out    vl_logic;
        wbLpEqexeSpAddr : out    vl_logic;
        exeMorMRpEqexeRpAddr: out    vl_logic;
        exeRTeqRA       : out    vl_logic;
        exeRTeqRB       : out    vl_logic;
        gprLpeqRp       : out    vl_logic;
        dcdRAL2         : in     vl_logic_vector(0 to 4);
        dcdRBL2         : in     vl_logic_vector(0 to 4);
        dcdRSRTL2       : in     vl_logic_vector(0 to 4);
        exeRS           : in     vl_logic_vector(0 to 4);
        exeApAddr       : in     vl_logic_vector(0 to 4);
        exeBpAddr       : in     vl_logic_vector(0 to 4);
        exeSpAddr       : in     vl_logic_vector(0 to 4);
        exeLpAddr       : in     vl_logic_vector(0 to 4);
        exeRpAddr       : in     vl_logic_vector(0 to 4);
        exeMacOrMultRpAddr: in     vl_logic_vector(0 to 4);
        wbLpAddr        : in     vl_logic_vector(0 to 4);
        PCL_wbRpAddr    : in     vl_logic_vector(0 to 4);
        PCL_lwbLpAddr   : in     vl_logic_vector(0 to 4);
        IFB_dcdFullL2   : in     vl_logic;
        exe1FullL2      : in     vl_logic;
        exe2FullL2      : in     vl_logic;
        wbFullL2        : in     vl_logic;
        lwbFullL2       : in     vl_logic;
        PCL_exeMacEnL2  : in     vl_logic;
        PCL_exeMultEnL2 : in     vl_logic;
        wbLpEqdcdSpAddr : out    vl_logic;
        lwbLpEqdcdSpAddr: out    vl_logic;
        exeMorMRpEqwbLpAddr: out    vl_logic;
        exeMorMRpEqlwbLpAddr: out    vl_logic;
        lwbLpAddr_NEG   : in     vl_logic_vector(0 to 4);
        wbRpAddr_NEG    : in     vl_logic_vector(0 to 4);
        sPortSelInc     : in     vl_logic;
        dcdBpMuxSel     : in     vl_logic;
        dcdSpMuxSel     : in     vl_logic;
        PCL_BpEqSp      : out    vl_logic
    );
end p405s_fileAddrCntl;
