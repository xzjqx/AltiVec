library verilog;
use verilog.vl_types.all;
entity p405s_mmu_utlb is
    port(
        DATA_COMP       : out    vl_logic;
        DO_00           : out    vl_logic;
        DO_01           : out    vl_logic;
        DO_02           : out    vl_logic;
        DO_03           : out    vl_logic;
        DO_04           : out    vl_logic;
        DO_05           : out    vl_logic;
        DO_06           : out    vl_logic;
        DO_07           : out    vl_logic;
        DO_08           : out    vl_logic;
        DO_09           : out    vl_logic;
        DO_10           : out    vl_logic;
        DO_11           : out    vl_logic;
        DO_12           : out    vl_logic;
        DO_13           : out    vl_logic;
        DO_14           : out    vl_logic;
        DO_15           : out    vl_logic;
        DO_16           : out    vl_logic;
        DO_17           : out    vl_logic;
        DO_18           : out    vl_logic;
        DO_19           : out    vl_logic;
        DO_20           : out    vl_logic;
        DO_21           : out    vl_logic;
        DO_E            : out    vl_logic;
        DO_G            : out    vl_logic;
        DO_I            : out    vl_logic;
        DO_K            : out    vl_logic;
        DO_M            : out    vl_logic;
        DO_PD_0         : out    vl_logic;
        DO_PD_1         : out    vl_logic;
        DO_PT_0         : out    vl_logic;
        DO_PT_1         : out    vl_logic;
        DO_PT_2         : out    vl_logic;
        DO_PT_3         : out    vl_logic;
        DO_V            : out    vl_logic;
        DO_W            : out    vl_logic;
        DSIZ_OUT_0      : out    vl_logic;
        DSIZ_OUT_1      : out    vl_logic;
        DSIZ_OUT_2      : out    vl_logic;
        DSIZ_OUT_3      : out    vl_logic;
        DSIZ_OUT_4      : out    vl_logic;
        DSIZ_OUT_5      : out    vl_logic;
        DSIZ_OUT_6      : out    vl_logic;
        DT_OUT          : out    vl_logic;
        EPN_OUT_00      : out    vl_logic;
        EPN_OUT_01      : out    vl_logic;
        EPN_OUT_02      : out    vl_logic;
        EPN_OUT_03      : out    vl_logic;
        EPN_OUT_04      : out    vl_logic;
        EPN_OUT_05      : out    vl_logic;
        EPN_OUT_06      : out    vl_logic;
        EPN_OUT_07      : out    vl_logic;
        EPN_OUT_08      : out    vl_logic;
        EPN_OUT_09      : out    vl_logic;
        EPN_OUT_10      : out    vl_logic;
        EPN_OUT_11      : out    vl_logic;
        EPN_OUT_12      : out    vl_logic;
        EPN_OUT_13      : out    vl_logic;
        EPN_OUT_14      : out    vl_logic;
        EPN_OUT_15      : out    vl_logic;
        EPN_OUT_16      : out    vl_logic;
        EPN_OUT_17      : out    vl_logic;
        EPN_OUT_18      : out    vl_logic;
        EPN_OUT_19      : out    vl_logic;
        EPN_OUT_20      : out    vl_logic;
        EPN_OUT_21      : out    vl_logic;
        EX_OUT          : out    vl_logic;
        INDEX_OUT_0     : out    vl_logic;
        INDEX_OUT_1     : out    vl_logic;
        INDEX_OUT_2     : out    vl_logic;
        INDEX_OUT_3     : out    vl_logic;
        INDEX_OUT_4     : out    vl_logic;
        INDEX_OUT_5     : out    vl_logic;
        MISS            : out    vl_logic;
        TAG_COMP        : out    vl_logic;
        TID_OUT_0       : out    vl_logic;
        TID_OUT_1       : out    vl_logic;
        TID_OUT_2       : out    vl_logic;
        TID_OUT_3       : out    vl_logic;
        TID_OUT_4       : out    vl_logic;
        TID_OUT_5       : out    vl_logic;
        TID_OUT_6       : out    vl_logic;
        TID_OUT_7       : out    vl_logic;
        WR_OUT          : out    vl_logic;
        ZSEL_OUT_0      : out    vl_logic;
        ZSEL_OUT_1      : out    vl_logic;
        ZSEL_OUT_2      : out    vl_logic;
        ZSEL_OUT_3      : out    vl_logic;
        DATA_EN         : in     vl_logic;
        DI_00           : in     vl_logic;
        DI_01           : in     vl_logic;
        DI_02           : in     vl_logic;
        DI_03           : in     vl_logic;
        DI_04           : in     vl_logic;
        DI_05           : in     vl_logic;
        DI_06           : in     vl_logic;
        DI_07           : in     vl_logic;
        DI_08           : in     vl_logic;
        DI_09           : in     vl_logic;
        DI_10           : in     vl_logic;
        DI_11           : in     vl_logic;
        DI_12           : in     vl_logic;
        DI_13           : in     vl_logic;
        DI_14           : in     vl_logic;
        DI_15           : in     vl_logic;
        DI_16           : in     vl_logic;
        DI_17           : in     vl_logic;
        DI_18           : in     vl_logic;
        DI_19           : in     vl_logic;
        DI_20           : in     vl_logic;
        DI_21           : in     vl_logic;
        DI_CI_00        : in     vl_logic;
        DI_CI_01        : in     vl_logic;
        DI_CI_02        : in     vl_logic;
        DI_CI_03        : in     vl_logic;
        DI_CI_04        : in     vl_logic;
        DI_CI_05        : in     vl_logic;
        DI_CI_06        : in     vl_logic;
        DI_CI_07        : in     vl_logic;
        DI_CI_08        : in     vl_logic;
        DI_CI_09        : in     vl_logic;
        DI_CI_10        : in     vl_logic;
        DI_CI_11        : in     vl_logic;
        DI_CI_12        : in     vl_logic;
        DI_CI_13        : in     vl_logic;
        DI_CI_14        : in     vl_logic;
        DI_CI_15        : in     vl_logic;
        DI_CI_16        : in     vl_logic;
        DI_CI_17        : in     vl_logic;
        DI_CI_18        : in     vl_logic;
        DI_CI_19        : in     vl_logic;
        DI_CI_20_TEST_EVEN: in     vl_logic;
        DI_CI_21_TEST_ODD: in     vl_logic;
        DI_E            : in     vl_logic;
        DI_G            : in     vl_logic;
        DI_I            : in     vl_logic;
        DI_K            : in     vl_logic;
        DI_M            : in     vl_logic;
        DI_PD_0         : in     vl_logic;
        DI_PD_1         : in     vl_logic;
        DI_PT_0         : in     vl_logic;
        DI_PT_1         : in     vl_logic;
        DI_PT_2         : in     vl_logic;
        DI_PT_3         : in     vl_logic;
        DI_V            : in     vl_logic;
        DI_W            : in     vl_logic;
        DSIZ_0          : in     vl_logic;
        DSIZ_1          : in     vl_logic;
        DSIZ_2          : in     vl_logic;
        DSIZ_3          : in     vl_logic;
        DSIZ_4          : in     vl_logic;
        DSIZ_5          : in     vl_logic;
        DSIZ_6          : in     vl_logic;
        DT              : in     vl_logic;
        DVS             : in     vl_logic;
        EN_ARRAYL1      : in     vl_logic;
        EN_C1           : in     vl_logic;
        EX              : in     vl_logic;
        INDEX_0         : in     vl_logic;
        INDEX_1         : in     vl_logic;
        INDEX_2         : in     vl_logic;
        INDEX_3         : in     vl_logic;
        INDEX_4         : in     vl_logic;
        INDEX_5         : in     vl_logic;
        INDEX_LOOKUPB   : in     vl_logic;
        INVAL           : in     vl_logic;
        RD_WRB          : in     vl_logic;
        SYS_CLK         : in     vl_logic;
        TAG_EN          : in     vl_logic;
        TEST_COMP       : in     vl_logic;
        TEST_M1         : in     vl_logic;
        TID_0           : in     vl_logic;
        TID_1           : in     vl_logic;
        TID_2           : in     vl_logic;
        TID_3           : in     vl_logic;
        TID_4           : in     vl_logic;
        TID_5           : in     vl_logic;
        TID_6           : in     vl_logic;
        TID_7           : in     vl_logic;
        WR              : in     vl_logic;
        ZSEL_0          : in     vl_logic;
        ZSEL_1          : in     vl_logic;
        ZSEL_2          : in     vl_logic;
        ZSEL_3          : in     vl_logic;
        reset           : in     vl_logic
    );
end p405s_mmu_utlb;
