library verilog;
use verilog.vl_types.all;
entity p405s_icu_PrControl is
    generic(
        iSideIdle       : integer := 2;
        iSideWa         : integer := 1;
        dSideIdle       : integer := 4;
        dSideLdCc       : integer := 2;
        dSideRd         : integer := 1;
        fillSmIdle      : integer := 32;
        fillSmReq       : integer := 16;
        fillSmFill      : integer := 8;
        fillSmWb        : integer := 4;
        fillSmWr0       : integer := 2;
        fillSmWr1       : integer := 1;
        preSmIdle       : integer := 16;
        preSmRd         : integer := 8;
        preSmWfr        : integer := 4;
        preSmReq        : integer := 2;
        preSmWf         : integer := 1;
        jtag0           : integer := 256;
        jtag1           : integer := 128;
        jtag2           : integer := 64;
        jtag3           : integer := 32;
        jtag4           : integer := 16;
        jtag5           : integer := 8;
        jtag6           : integer := 4;
        jtag7           : integer := 2;
        jtag8           : integer := 1
    );
    port(
        ICU_request_NEG : out    vl_logic;
        ICU_size_NEG    : out    vl_logic_vector(0 to 1);
        ICU_Abort_NEG   : out    vl_logic;
        ICU_cacheable_NEG: out    vl_logic;
        ICU_ocmReqPending_NEG: out    vl_logic;
        ICU_isCA        : out    vl_logic;
        ICU_dsCA        : out    vl_logic;
        ICU_sleepReq    : out    vl_logic;
        ICU_syncAfterReset: out    vl_logic;
        ICU_ifbError    : out    vl_logic_vector(0 to 1);
        ICU_mmuRdarE2   : out    vl_logic;
        tagVSel_1       : out    vl_logic;
        lruRdSel        : out    vl_logic;
        dataCcSel       : out    vl_logic_vector(0 to 3);
        plbLowSel       : out    vl_logic_vector(0 to 1);
        plbHighSel      : out    vl_logic_vector(0 to 1);
        rarsSel         : out    vl_logic_vector(0 to 1);
        vcarsSel        : out    vl_logic_vector(0 to 1);
        dsRdMuxSel      : out    vl_logic;
        vcarE2          : out    vl_logic;
        isU0AttrL2      : out    vl_logic;
        cdbdrE1         : out    vl_logic;
        fillWr0L2       : out    vl_logic;
        vcarsCCE2       : out    vl_logic;
        vcarInSelL2     : out    vl_logic;
        vcarspSel       : out    vl_logic_vector(0 to 1);
        icuRdarE1       : out    vl_logic;
        icuRdarE2       : out    vl_logic;
        dsVcar1E2       : out    vl_logic;
        dsVcar2E2       : out    vl_logic;
        isBusSel        : out    vl_logic_vector(0 to 1);
        Lx27Sel         : out    vl_logic;
        Lx28Sel         : out    vl_logic;
        Lx29Sel         : out    vl_logic;
        lruRdCcE1       : out    vl_logic;
        VaVbWrE1        : out    vl_logic;
        vcarSel_pri_NEG : in     vl_logic;
        tagBWE1         : out    vl_logic;
        wbHighE2        : out    vl_logic_vector(0 to 3);
        wbLowE2         : out    vl_logic;
        wbTagE1         : out    vl_logic;
        fillAE2         : out    vl_logic_vector(0 to 7);
        fillBE2         : out    vl_logic_vector(0 to 7);
        newLruBitIn     : out    vl_logic;
        wrVaIn          : out    vl_logic;
        newVaBitIn      : out    vl_logic;
        wrVbIn          : out    vl_logic;
        newVbBitIn      : out    vl_logic;
        dataRdWrRegIn   : out    vl_logic;
        tagRdWrRegIn    : out    vl_logic;
        wrATagNotB      : out    vl_logic;
        vaOutL2         : out    vl_logic;
        vbOutL2         : out    vl_logic;
        eo_y_NEG        : out    vl_logic;
        eo_z_NEG        : out    vl_logic;
        eo_r            : out    vl_logic;
        eo_q            : out    vl_logic;
        rdStateL2       : out    vl_logic;
        dsRD1cycle      : out    vl_logic;
        wrFlashIn       : out    vl_logic;
        resetCore2L2    : out    vl_logic;
        sc3L2           : out    vl_logic;
        jtag2ndWr       : out    vl_logic;
        diagBus         : out    vl_logic_vector(0 to 22);
        rdOrWaAndXltValid: out    vl_logic;
        frAndDsRdy      : out    vl_logic;
        cycle_RA_p3_NEG : out    vl_logic;
        cycle_RB_p3_NEG : out    vl_logic;
        cycle_RT_p3_NEG : out    vl_logic;
        cycle_parity_p3_NEG: out    vl_logic;
        forceNlL2       : out    vl_logic;
        setForceNl      : out    vl_logic;
        rdSt_RDA_pg4_NEG: out    vl_logic;
        VaVb_VR_pg4_NEG : out    vl_logic;
        bufValidL2_NEG  : out    vl_logic;
        ldcc2RdNoAb_NEG : out    vl_logic;
        wrLruNoHit_NEG  : out    vl_logic;
        nfr_ABC_p2_NEG  : out    vl_logic;
        eo_z2_NEG       : out    vl_logic;
        lxFetchValidIn_A_NEG: out    vl_logic;
        lxFetchValidIn_B_NEG: out    vl_logic;
        lxSel_C_NEG     : out    vl_logic;
        lxSel_D_NEG     : out    vl_logic;
        lxFetchValidL2  : out    vl_logic;
        vcarSel_noEO    : out    vl_logic;
        tagSelBit0_E_NEG: out    vl_logic;
        tagSelBit0_F_NEG: out    vl_logic;
        ocmDvQ_1_NEG    : out    vl_logic;
        nxtWa_W_NEG     : out    vl_logic;
        nxtWa_X_NEG     : out    vl_logic;
        missL2          : out    vl_logic;
        PCL_mtSPR       : in     vl_logic;
        PLB_icuAddrAck  : in     vl_logic;
        PLB_icuRdDAck   : in     vl_logic;
        PLB_icuError    : in     vl_logic;
        PLB_icuBusy     : in     vl_logic;
        PLB_dcuBusy     : in     vl_logic;
        PLB_icuRdWrAddr : in     vl_logic_vector(1 to 3);
        PLB_sSize       : in     vl_logic;
        PLB_sampleCycle : in     vl_logic;
        OCM_isDValid    : in     vl_logic_vector(0 to 1);
        OCM_isHold      : in     vl_logic;
        IFB_fetchReq    : in     vl_logic;
        df_cpuEa        : in     vl_logic_vector(27 to 29);
        IFB_isNL        : in     vl_logic;
        IFB_isAbort     : in     vl_logic_vector(0 to 2);
        IFB_icuCancelData: in     vl_logic;
        PCL_icuOp       : in     vl_logic_vector(0 to 3);
        VCT_icuWbAbort  : in     vl_logic;
        VCT_exeAbort    : in     vl_logic;
        IFB_cntxSync    : in     vl_logic;
        MMU_isDsXltValidL2: in     vl_logic;
        MMU_isDsCacheableL2: in     vl_logic;
        MMU_icuDsAbort  : in     vl_logic;
        MMU_isXltValid_NEG: in     vl_logic;
        MMU_isCacheable : in     vl_logic_vector(1 to 2);
        MMU_icuIsAbort  : in     vl_logic;
        MMU_isU0Attr    : in     vl_logic;
        df_preFetchEnable: in     vl_logic;
        df_forceOnly1Req: in     vl_logic;
        df_ftchMissBlkWr: in     vl_logic;
        df_nonC_8       : in     vl_logic;
        df_nonCpreFetchEn: in     vl_logic;
        df_plbaOverflow : in     vl_logic;
        df_vcarVcarsCompare: in     vl_logic;
        df_plb27L2      : in     vl_logic;
        compB_NEG       : in     vl_logic;
        compAlru_NEG    : in     vl_logic;
        dsCompA         : in     vl_logic;
        dsCompB         : in     vl_logic;
        lruOut          : in     vl_logic;
        vaOut           : in     vl_logic;
        vbOut           : in     vl_logic;
        forceNlIn       : in     vl_logic;
        rdStateIn       : in     vl_logic;
        nxtFetchRd      : in     vl_logic;
        lxSel           : in     vl_logic;
        lxFetchValidIn  : in     vl_logic;
        nxtWait         : in     vl_logic;
        bufValidIn_NEG  : in     vl_logic;
        df_selCCR0      : in     vl_logic;
        JTG_iCacheWr    : in     vl_logic;
        icuTagDataSel   : in     vl_logic;
        icuBaSel        : in     vl_logic;
        CB              : in     vl_logic;
        resetCoreIn     : in     vl_logic;
        testEn_NEG      : in     vl_logic;
        missIn          : in     vl_logic;
        PLB_sampleCycleAlt: in     vl_logic;
        CPM_c405SyncBypass: in     vl_logic
    );
end p405s_icu_PrControl;
