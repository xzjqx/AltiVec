library verilog;
use verilog.vl_types.all;
entity PPC405F5V1_soft is
    port(
        C405_apuDcdFull : out    vl_logic;
        C405_apuDcdHold : out    vl_logic;
        C405_apuDcdInstruction: out    vl_logic_vector(0 to 31);
        C405_apuExeFlush: out    vl_logic;
        C405_apuExeHold : out    vl_logic;
        C405_apuExeLoadDBus: out    vl_logic_vector(0 to 31);
        C405_apuExeLoadDValid: out    vl_logic;
        C405_apuExeRaData: out    vl_logic_vector(0 to 31);
        C405_apuExeRbData: out    vl_logic_vector(0 to 31);
        C405_apuExeWdCnt: out    vl_logic_vector(0 to 1);
        C405_apuMsrFE0  : out    vl_logic;
        C405_apuMsrFE1  : out    vl_logic;
        C405_apuWbByteEn: out    vl_logic_vector(0 to 3);
        C405_apuWbEndian: out    vl_logic;
        C405_apuWbFlush : out    vl_logic;
        C405_apuWbHold  : out    vl_logic;
        C405_apuXerCA   : out    vl_logic;
        C405_cpmCoreSleepReq: out    vl_logic;
        C405_cpmMsrCE   : out    vl_logic;
        C405_cpmMsrEE   : out    vl_logic;
        C405_cpmTimerIRQ: out    vl_logic;
        C405_cpmTimerResetReq: out    vl_logic;
        C405_dbgLoadDataOnApuDBus: out    vl_logic;
        C405_dbgMsrWE   : out    vl_logic;
        C405_dbgStopAck : out    vl_logic;
        C405_dbgWbComplete: out    vl_logic;
        C405_dbgWbFull  : out    vl_logic;
        C405_dbgWbIar   : out    vl_logic_vector(0 to 29);
        C405_dcrABus    : out    vl_logic_vector(0 to 9);
        C405_dcrDBusOut : out    vl_logic_vector(0 to 31);
        C405_dcrRead    : out    vl_logic;
        C405_dcrWrite   : out    vl_logic;
        C405_dsocmAbortOp: out    vl_logic;
        C405_dsocmAbortReq: out    vl_logic;
        C405_dsocmABus  : out    vl_logic_vector(0 to 29);
        C405_dsocmByteEn: out    vl_logic_vector(0 to 3);
        C405_dsocmCacheable: out    vl_logic;
        C405_dsocmGuarded: out    vl_logic;
        C405_dsocmLoadReq: out    vl_logic;
        C405_dsocmStoreReq: out    vl_logic;
        C405_dsocmStringMultiple: out    vl_logic;
        C405_dsocmU0Attr: out    vl_logic;
        C405_dsocmWait  : out    vl_logic;
        C405_dsocmWrDBus: out    vl_logic_vector(0 to 31);
        C405_dsocmXlateValid: out    vl_logic;
        C405_isocmAbort : out    vl_logic;
        C405_isocmABus  : out    vl_logic_vector(0 to 29);
        C405_isocmCacheable: out    vl_logic;
        C405_isocmContextSync: out    vl_logic;
        C405_isocmIcuReady: out    vl_logic;
        C405_isocmReqPending: out    vl_logic;
        C405_isocmU0Attr: out    vl_logic;
        C405_isocmXlateValid: out    vl_logic;
        C405_jtgCaptureDR: out    vl_logic;
        C405_jtgExtest  : out    vl_logic;
        C405_jtgPgmOut  : out    vl_logic;
        C405_jtgShiftDR : out    vl_logic;
        C405_jtgTDO     : out    vl_logic;
        C405_jtgTDOEn   : out    vl_logic;
        C405_jtgUpdateDR: out    vl_logic;
        C405_testDiagAbistDone: out    vl_logic;
        C405_testScanOut: out    vl_logic_vector(0 to 7);
        C405_plbDcuAbort: out    vl_logic;
        C405_plbDcuABus : out    vl_logic_vector(0 to 31);
        C405_plbDcuBE   : out    vl_logic_vector(0 to 7);
        C405_plbDcuCacheable: out    vl_logic;
        C405_plbDcuGuarded: out    vl_logic;
        C405_plbDcuPriority: out    vl_logic_vector(0 to 1);
        C405_plbDcuRequest: out    vl_logic;
        C405_plbDcuRNW  : out    vl_logic;
        C405_plbDcuSize2: out    vl_logic;
        C405_plbDcuU0Attr: out    vl_logic;
        C405_plbDcuWrDBus: out    vl_logic_vector(0 to 63);
        C405_plbDcuWriteThru: out    vl_logic;
        C405_plbIcuAbort: out    vl_logic;
        C405_plbIcuABus : out    vl_logic_vector(0 to 29);
        C405_plbIcuCacheable: out    vl_logic;
        C405_plbIcuPriority: out    vl_logic_vector(0 to 1);
        C405_plbIcuRequest: out    vl_logic;
        C405_plbIcuSize : out    vl_logic_vector(2 to 3);
        C405_plbIcuU0Attr: out    vl_logic;
        C405_rstChipResetReq: out    vl_logic;
        C405_rstCoreResetReq: out    vl_logic;
        C405_rstSystemResetReq: out    vl_logic;
        C405_trcCycle   : out    vl_logic;
        C405_trcEvenExecutionStatus: out    vl_logic_vector(0 to 1);
        C405_trcOddExecutionStatus: out    vl_logic_vector(0 to 1);
        C405_trcTraceStatus: out    vl_logic_vector(0 to 3);
        C405_trcTriggerEventOut: out    vl_logic;
        C405_trcTriggerEventType: out    vl_logic_vector(0 to 10);
        C405_xxxMachineCheck: out    vl_logic;
        APU_c405DcdApuOp: in     vl_logic;
        APU_c405DcdCREn : in     vl_logic;
        APU_c405DcdForceAlgn: in     vl_logic;
        APU_c405DcdForceBESteering: in     vl_logic;
        APU_c405DcdFpuOp: in     vl_logic;
        APU_c405DcdGprWrite: in     vl_logic;
        APU_c405DcdLdStByte: in     vl_logic;
        APU_c405DcdLdStDw: in     vl_logic;
        APU_c405DcdLdStHw: in     vl_logic;
        APU_c405DcdLdStQw: in     vl_logic;
        APU_c405DcdLdStWd: in     vl_logic;
        APU_c405DcdLoad : in     vl_logic;
        APU_c405DcdPrivOp: in     vl_logic;
        APU_c405DcdRaEn : in     vl_logic;
        APU_c405DcdRbEn : in     vl_logic;
        APU_c405DcdStore: in     vl_logic;
        APU_c405DcdTrapBE: in     vl_logic;
        APU_c405DcdTrapLE: in     vl_logic;
        APU_c405DcdUpdate: in     vl_logic;
        APU_c405DcdValidOp: in     vl_logic;
        APU_c405DcdXerCAEn: in     vl_logic;
        APU_c405DcdXerOVEn: in     vl_logic;
        APU_c405Exception: in     vl_logic;
        APU_c405ExeBlockingMCO: in     vl_logic;
        APU_c405ExeBusy : in     vl_logic;
        APU_c405ExeCR   : in     vl_logic_vector(0 to 3);
        APU_c405ExeCRField: in     vl_logic_vector(0 to 2);
        APU_c405ExeLdDepend: in     vl_logic;
        APU_c405ExeNonBlockingMCO: in     vl_logic;
        APU_c405ExeResult: in     vl_logic_vector(0 to 31);
        APU_c405ExeXerCA: in     vl_logic;
        APU_c405ExeXerOV: in     vl_logic;
        APU_c405FpuException: in     vl_logic;
        APU_c405LwbLdDepend: in     vl_logic;
        APU_c405SleepReq: in     vl_logic;
        APU_c405WbLdDepend: in     vl_logic;
        CPM_c405Clock   : in     vl_logic;
        CPM_c405CoreClkInactive: in     vl_logic;
        CPM_c405CpuClkEn_CClk: in     vl_logic;
        CPM_c405JtagClkEn_CClk: in     vl_logic;
        CPM_c405PlbSampleCycle: in     vl_logic;
        CPM_c405PlbSampleCycleAlt: in     vl_logic;
        CPM_c405PlbSyncClock: in     vl_logic;
        CPM_c405SyncBypass: in     vl_logic;
        CPM_c405TimerClkEn_CClk: in     vl_logic;
        CPM_c405TimerTick: in     vl_logic;
        DBG_c405DebugHalt: in     vl_logic;
        DBG_c405ExtBusHoldAck: in     vl_logic;
        DBG_c405UncondDebugEvent: in     vl_logic;
        DCR_c405Ack     : in     vl_logic;
        DCR_c405DBusIn  : in     vl_logic_vector(0 to 31);
        DSOCM_c405Complete: in     vl_logic;
        DSOCM_c405DisOperandFwd: in     vl_logic;
        DSOCM_c405Hold  : in     vl_logic;
        DSOCM_c405RdDBus: in     vl_logic_vector(0 to 31);
        EIC_c405CritInputIRQ: in     vl_logic;
        EIC_c405ExtInputIRQ: in     vl_logic;
        ISOCM_c405Hold  : in     vl_logic;
        ISOCM_c405RdDBus: in     vl_logic_vector(0 to 63);
        ISOCM_c405RdDValid: in     vl_logic_vector(0 to 1);
        JTG_c405BndScanTDO: in     vl_logic;
        JTG_c405TCK     : in     vl_logic;
        JTG_c405TDI     : in     vl_logic;
        JTG_c405TMS     : in     vl_logic;
        JTG_c405TRST_NEG: in     vl_logic;
        TEST_c405BistCClk: in     vl_logic;
        TEST_c405BistCE0StClk: in     vl_logic;
        TEST_c405BistCE1Enable: in     vl_logic;
        TEST_c405BistCE1Mode: in     vl_logic;
        TEST_c405CE0EVS : in     vl_logic;
        TEST_c405CntlPoint: in     vl_logic;
        TEST_c405ScanEnable: in     vl_logic;
        TEST_c405ScanIn : in     vl_logic_vector(0 to 7);
        TEST_c405TestM1 : in     vl_logic;
        TEST_c405TestM3 : in     vl_logic;
        TEST_c405TestMode: in     vl_logic;
        PLB_c405DcuAddrAck: in     vl_logic;
        PLB_c405DcuBusy : in     vl_logic;
        PLB_c405DcuErr  : in     vl_logic;
        PLB_c405DcuRdDAck: in     vl_logic;
        PLB_c405DcuRdDBus: in     vl_logic_vector(0 to 63);
        PLB_c405DcuRdWdAddr: in     vl_logic_vector(1 to 3);
        PLB_c405DcuSSize1: in     vl_logic;
        PLB_c405DcuWrDAck: in     vl_logic;
        PLB_c405IcuAddrAck: in     vl_logic;
        PLB_c405IcuBusy : in     vl_logic;
        PLB_c405IcuErr  : in     vl_logic;
        PLB_c405IcuRdDAck: in     vl_logic;
        PLB_c405IcuRdDBus: in     vl_logic_vector(0 to 63);
        PLB_c405IcuRdWdAddr: in     vl_logic_vector(1 to 3);
        PLB_c405IcuSSize1: in     vl_logic;
        RST_c405ResetChip: in     vl_logic;
        RST_c405ResetCore: in     vl_logic;
        RST_c405ResetSystem: in     vl_logic;
        TIE_c405ApuDivEn: in     vl_logic;
        TIE_c405ApuPresent: in     vl_logic;
        TIE_c405ClockEnable: in     vl_logic;
        TIE_c405DeterministicMult: in     vl_logic;
        TIE_c405DisOperandFwd: in     vl_logic;
        TIE_c405DutyEnable: in     vl_logic;
        TIE_c405MmuEn   : in     vl_logic;
        TIE_c405PVR     : in     vl_logic_vector(0 to 31);
        TRC_c405TraceDisable: in     vl_logic;
        TRC_c405TriggerEventIn: in     vl_logic;
        C405_bistPepsPF : out    vl_logic_vector(0 to 2);
        BIST_c405dcuBistDebugEn: in     vl_logic_vector(3 downto 0);
        BIST_c405dcuBistDebugSi: in     vl_logic_vector(3 downto 0);
        BIST_c405dcuBistMbRun: in     vl_logic;
        BIST_c405dcuBistModeRegIn: in     vl_logic_vector(18 downto 0);
        BIST_c405dcuBistModeRegSi: in     vl_logic;
        BIST_c405dcuBistParallelDr: in     vl_logic;
        BIST_c405dcuBistShiftDr: in     vl_logic;
        BIST_c405icuBistDebugEn: in     vl_logic_vector(3 downto 0);
        BIST_c405icuBistDebugSi: in     vl_logic_vector(3 downto 0);
        BIST_c405icuBistMbRun: in     vl_logic;
        BIST_c405icuBistModeRegIn: in     vl_logic_vector(18 downto 0);
        BIST_c405icuBistModeRegSi: in     vl_logic;
        BIST_c405icuBistParallelDr: in     vl_logic;
        BIST_c405icuBistShiftDr: in     vl_logic;
        C405_bistdcuBistDebugSo: out    vl_logic_vector(3 downto 0);
        C405_bistdcuBistModeRegSo: out    vl_logic;
        C405_bistdcuBistModeRegOut: out    vl_logic_vector(18 downto 0);
        C405_bisticuBistDebugSo: out    vl_logic_vector(3 downto 0);
        C405_bisticuBistModeRegSo: out    vl_logic;
        C405_bisticuBistModeRegOut: out    vl_logic_vector(18 downto 0)
    );
end PPC405F5V1_soft;
