// 
// ************************************************************************** 
// 
//  Copyright (c) International Business Machines Corporation, 2005. 
// 
//  This file contains trade secrets and other proprietary and confidential 
//  information of International Business Machines Corporation which are 
//  protected by copyright and other intellectual property rights and shall 
//  not be reproduced, transferred to other documents, disclosed to others, 
//  or used for any purpose except as specifically authorized in writing by 
//  International Business Machines Corporation. This notice must be 
//  contained as part of this text at all times. 
// 
// ************************************************************************** 
//
module PPC405F5V1_soft( C405_apuDcdFull, C405_apuDcdHold, C405_apuDcdInstruction,
     C405_apuExeFlush, C405_apuExeHold, C405_apuExeLoadDBus, C405_apuExeLoadDValid,
     C405_apuExeRaData, C405_apuExeRbData, C405_apuExeWdCnt, C405_apuMsrFE0,
     C405_apuMsrFE1, C405_apuWbByteEn, C405_apuWbEndian, C405_apuWbFlush, C405_apuWbHold,
     C405_apuXerCA, C405_cpmCoreSleepReq, C405_cpmMsrCE, C405_cpmMsrEE, C405_cpmTimerIRQ,
     C405_cpmTimerResetReq, C405_dbgLoadDataOnApuDBus, C405_dbgMsrWE, C405_dbgStopAck,
     C405_dbgWbComplete, C405_dbgWbFull, C405_dbgWbIar, C405_dcrABus,
     C405_dcrDBusOut, C405_dcrRead, C405_dcrWrite, 
     C405_dsocmAbortOp, C405_dsocmAbortReq,C405_dsocmABus, C405_dsocmByteEn, C405_dsocmCacheable,
     C405_dsocmGuarded, C405_dsocmLoadReq, C405_dsocmStoreReq, C405_dsocmStringMultiple,
     C405_dsocmU0Attr, C405_dsocmWait, C405_dsocmWrDBus, C405_dsocmXlateValid,
      C405_isocmAbort,C405_isocmABus, C405_isocmCacheable, C405_isocmContextSync,
     C405_isocmIcuReady, C405_isocmReqPending, C405_isocmU0Attr, C405_isocmXlateValid,
     C405_jtgCaptureDR, C405_jtgExtest, C405_jtgPgmOut, C405_jtgShiftDR, C405_jtgTDO,
     C405_jtgTDOEn, C405_jtgUpdateDR, C405_testDiagAbistDone, 
     C405_testScanOut, C405_plbDcuAbort,C405_plbDcuABus,  C405_plbDcuBE,
     C405_plbDcuCacheable, C405_plbDcuGuarded, C405_plbDcuPriority, C405_plbDcuRequest,
	 C405_plbDcuRNW,C405_plbDcuSize2, C405_plbDcuU0Attr, C405_plbDcuWrDBus,
     C405_plbDcuWriteThru, C405_plbIcuAbort,C405_plbIcuABus,  C405_plbIcuCacheable,
     C405_plbIcuPriority, C405_plbIcuRequest, C405_plbIcuSize, C405_plbIcuU0Attr,
     C405_rstChipResetReq, C405_rstCoreResetReq, C405_rstSystemResetReq, C405_trcCycle,
     C405_trcEvenExecutionStatus, C405_trcOddExecutionStatus,
     C405_trcTraceStatus, C405_trcTriggerEventOut, C405_trcTriggerEventType,
     C405_xxxMachineCheck,
     APU_c405DcdApuOp, APU_c405DcdCREn, APU_c405DcdForceAlgn,
     APU_c405DcdForceBESteering, APU_c405DcdFpuOp, APU_c405DcdGprWrite, APU_c405DcdLdStByte,
     APU_c405DcdLdStDw, APU_c405DcdLdStHw, APU_c405DcdLdStQw, APU_c405DcdLdStWd,
     APU_c405DcdLoad, APU_c405DcdPrivOp, APU_c405DcdRaEn, APU_c405DcdRbEn, APU_c405DcdStore,
     APU_c405DcdTrapBE, APU_c405DcdTrapLE, APU_c405DcdUpdate, APU_c405DcdValidOp,
     APU_c405DcdXerCAEn, APU_c405DcdXerOVEn, APU_c405Exception, APU_c405ExeBlockingMCO,
     APU_c405ExeBusy, APU_c405ExeCR, APU_c405ExeCRField, APU_c405ExeLdDepend,
     APU_c405ExeNonBlockingMCO, APU_c405ExeResult, APU_c405ExeXerCA, APU_c405ExeXerOV,
     APU_c405FpuException, APU_c405LwbLdDepend, APU_c405SleepReq, APU_c405WbLdDepend,
     CPM_c405Clock, CPM_c405CoreClkInactive,CPM_c405CpuClkEn_CClk,CPM_c405JtagClkEn_CClk,
     CPM_c405PlbSampleCycle,CPM_c405PlbSampleCycleAlt,CPM_c405PlbSyncClock,CPM_c405SyncBypass,
	 CPM_c405TimerClkEn_CClk,CPM_c405TimerTick, 
	 DBG_c405DebugHalt, DBG_c405ExtBusHoldAck, DBG_c405UncondDebugEvent,
     DCR_c405Ack, DCR_c405DBusIn, DSOCM_c405Complete, DSOCM_c405DisOperandFwd,
     DSOCM_c405Hold, DSOCM_c405RdDBus, EIC_c405CritInputIRQ, EIC_c405ExtInputIRQ,
     ISOCM_c405Hold, ISOCM_c405RdDBus, ISOCM_c405RdDValid, JTG_c405BndScanTDO,
     JTG_c405TCK, JTG_c405TDI, JTG_c405TMS, JTG_c405TRST_NEG,
     TEST_c405BistCClk,TEST_c405BistCE0StClk,TEST_c405BistCE1Enable,TEST_c405BistCE1Mode,
	 TEST_c405CE0EVS,TEST_c405CntlPoint,TEST_c405ScanEnable,TEST_c405ScanIn, 
	  TEST_c405TestM1, TEST_c405TestM3,TEST_c405TestMode,
     PLB_c405DcuAddrAck, PLB_c405DcuBusy, PLB_c405DcuErr, PLB_c405DcuRdDAck,
     PLB_c405DcuRdDBus, PLB_c405DcuRdWdAddr, PLB_c405DcuSSize1, PLB_c405DcuWrDAck,
     PLB_c405IcuAddrAck, PLB_c405IcuBusy, PLB_c405IcuErr, PLB_c405IcuRdDAck,
     PLB_c405IcuRdDBus, PLB_c405IcuRdWdAddr, PLB_c405IcuSSize1, RST_c405ResetChip,
     RST_c405ResetCore, RST_c405ResetSystem, TIE_c405ApuDivEn, TIE_c405ApuPresent,
     TIE_c405ClockEnable,TIE_c405DeterministicMult, TIE_c405DisOperandFwd,TIE_c405DutyEnable,
	 TIE_c405MmuEn, TIE_c405PVR,TRC_c405TraceDisable, TRC_c405TriggerEventIn, 
	 C405_bistPepsPF,
	 BIST_c405dcuBistDebugEn,
	 BIST_c405dcuBistDebugSi,
     BIST_c405dcuBistMbRun,
     BIST_c405dcuBistModeRegIn,
     BIST_c405dcuBistModeRegSi,
	 BIST_c405dcuBistParallelDr,
	 BIST_c405dcuBistShiftDr,
	 BIST_c405icuBistDebugEn,
	 BIST_c405icuBistDebugSi,
	 BIST_c405icuBistMbRun,
	 BIST_c405icuBistModeRegIn,
	 BIST_c405icuBistModeRegSi,
	 BIST_c405icuBistParallelDr,
	 BIST_c405icuBistShiftDr,
     C405_bistdcuBistDebugSo,
     C405_bistdcuBistModeRegSo,
     C405_bistdcuBistModeRegOut,
     C405_bisticuBistDebugSo,        
     C405_bisticuBistModeRegSo,   
     C405_bisticuBistModeRegOut );


output  C405_apuDcdFull, C405_apuDcdHold, C405_apuExeFlush, C405_apuExeHold,
     C405_apuExeLoadDValid, C405_apuMsrFE0, C405_apuMsrFE1, C405_apuWbEndian, C405_apuWbFlush,
     C405_apuWbHold, C405_apuXerCA, C405_cpmCoreSleepReq, C405_cpmMsrCE, C405_cpmMsrEE,
     C405_cpmTimerIRQ, C405_cpmTimerResetReq, C405_dbgLoadDataOnApuDBus, C405_dbgMsrWE,
     C405_dbgStopAck, C405_dbgWbComplete, C405_dbgWbFull, C405_dcrRead, C405_dcrWrite,
     C405_dsocmAbortOp, C405_dsocmAbortReq, C405_dsocmCacheable, C405_dsocmGuarded,
     C405_dsocmLoadReq, C405_dsocmStoreReq, C405_dsocmStringMultiple, C405_dsocmU0Attr,
     C405_dsocmWait, C405_dsocmXlateValid, C405_isocmAbort, C405_isocmCacheable,
     C405_isocmContextSync, C405_isocmIcuReady, C405_isocmReqPending, C405_isocmU0Attr,
     C405_isocmXlateValid, C405_jtgCaptureDR, C405_jtgExtest, C405_jtgPgmOut, C405_jtgShiftDR,
     C405_jtgTDO, C405_jtgTDOEn, C405_jtgUpdateDR, C405_testDiagAbistDone, 
     C405_plbDcuAbort, C405_plbDcuCacheable, C405_plbDcuGuarded, C405_plbDcuRNW,
     C405_plbDcuRequest, C405_plbDcuSize2, C405_plbDcuU0Attr, C405_plbDcuWriteThru,
     C405_plbIcuAbort, C405_plbIcuCacheable, C405_plbIcuRequest, C405_plbIcuU0Attr,
     C405_rstChipResetReq, C405_rstCoreResetReq, C405_rstSystemResetReq, C405_trcCycle,
     C405_trcTriggerEventOut, C405_xxxMachineCheck;


input  APU_c405DcdApuOp, APU_c405DcdCREn, APU_c405DcdForceAlgn, APU_c405DcdForceBESteering,
     APU_c405DcdFpuOp, APU_c405DcdGprWrite, APU_c405DcdLdStByte, APU_c405DcdLdStDw,
     APU_c405DcdLdStHw, APU_c405DcdLdStQw, APU_c405DcdLdStWd, APU_c405DcdLoad,
     APU_c405DcdPrivOp, APU_c405DcdRaEn, APU_c405DcdRbEn, APU_c405DcdStore, APU_c405DcdTrapBE,
     APU_c405DcdTrapLE, APU_c405DcdUpdate, APU_c405DcdValidOp, APU_c405DcdXerCAEn,
     APU_c405DcdXerOVEn, APU_c405Exception, APU_c405ExeBlockingMCO, APU_c405ExeBusy,
	 
     APU_c405ExeLdDepend, APU_c405ExeNonBlockingMCO, APU_c405ExeXerCA, APU_c405ExeXerOV,
     APU_c405FpuException, APU_c405LwbLdDepend, APU_c405SleepReq, APU_c405WbLdDepend,
     CPM_c405Clock, CPM_c405CoreClkInactive,CPM_c405CpuClkEn_CClk,CPM_c405JtagClkEn_CClk,
     CPM_c405PlbSampleCycle,CPM_c405TimerClkEn_CClk,
     CPM_c405TimerTick, DBG_c405DebugHalt, DBG_c405ExtBusHoldAck, DBG_c405UncondDebugEvent,
     DCR_c405Ack, DSOCM_c405Complete, DSOCM_c405DisOperandFwd, DSOCM_c405Hold,
     EIC_c405CritInputIRQ, EIC_c405ExtInputIRQ, ISOCM_c405Hold, JTG_c405BndScanTDO,
     JTG_c405TCK, JTG_c405TDI, JTG_c405TMS, JTG_c405TRST_NEG,
     TEST_c405BistCClk,
     TEST_c405CntlPoint, TEST_c405TestM1, TEST_c405TestM3, PLB_c405DcuAddrAck, PLB_c405DcuBusy,
     PLB_c405DcuErr, PLB_c405DcuRdDAck, PLB_c405DcuSSize1, PLB_c405DcuWrDAck,
     PLB_c405IcuAddrAck, PLB_c405IcuBusy, PLB_c405IcuErr, PLB_c405IcuRdDAck, PLB_c405IcuSSize1,
     RST_c405ResetChip, RST_c405ResetCore, RST_c405ResetSystem, TIE_c405ApuDivEn,
     TIE_c405ApuPresent, TIE_c405DeterministicMult, TIE_c405DisOperandFwd, TIE_c405MmuEn,
     TRC_c405TraceDisable, TRC_c405TriggerEventIn, TEST_c405CE0EVS,  
     TEST_c405BistCE0StClk, TEST_c405BistCE1Enable, TEST_c405BistCE1Mode,
     TIE_c405ClockEnable, TIE_c405DutyEnable;

// added for tbird
input          CPM_c405SyncBypass;
input          CPM_c405PlbSyncClock;
input          CPM_c405PlbSampleCycleAlt;
 
output [0:31]  C405_apuDcdInstruction;
output [0:29]  C405_dsocmABus;
output [0:31]  C405_dcrDBusOut;
output [0:31]  C405_apuExeRbData;
output [0:31]  C405_apuExeLoadDBus;
output [0:3]  C405_apuWbByteEn;
output [0:1]  C405_plbDcuPriority;
output [0:1]  C405_trcOddExecutionStatus;
output [0:10]  C405_trcTriggerEventType;
output [0:7]  C405_plbDcuBE;
output [0:63]  C405_plbDcuWrDBus;
output [0:31]  C405_plbDcuABus;
output [2:3]  C405_plbIcuSize;
output [0:29]  C405_plbIcuABus;
output [0:7]  C405_testScanOut;
output [0:3]  C405_dsocmByteEn;
output [0:29]  C405_isocmABus;
output [0:1]  C405_plbIcuPriority;
output [0:31]  C405_dsocmWrDBus;
output [0:3]  C405_trcTraceStatus;
output [0:1]  C405_trcEvenExecutionStatus;
output [0:29]  C405_dbgWbIar;
output [0:9]  C405_dcrABus;
output [0:1]  C405_apuExeWdCnt;
output [0:31]  C405_apuExeRaData;
output [0:2]  C405_bistPepsPF;

input [0:31]  DSOCM_c405RdDBus;
input [0:3]  APU_c405ExeCR;
input [0:63]  ISOCM_c405RdDBus;
input [0:31]  APU_c405ExeResult;
input [0:2]  APU_c405ExeCRField;
input [0:31]  TIE_c405PVR;
input [1:3]  PLB_c405DcuRdWdAddr;
input [0:63]  PLB_c405DcuRdDBus;
input [0:31]  DCR_c405DBusIn;
input [1:3]  PLB_c405IcuRdWdAddr;
input [0:63]  PLB_c405IcuRdDBus;
input [0:1]  ISOCM_c405RdDValid;
input [0:7]  TEST_c405ScanIn;
input   TEST_c405ScanEnable;
input   TEST_c405TestMode;


// Bist Interface
input          BIST_c405dcuBistMbRun;

input  [3:0]   BIST_c405dcuBistDebugSi;
input  [3:0]   BIST_c405dcuBistDebugEn;
output [3:0]   C405_bistdcuBistDebugSo;

input          BIST_c405dcuBistShiftDr;
input          BIST_c405dcuBistModeRegSi;
output         C405_bistdcuBistModeRegSo;

input          BIST_c405dcuBistParallelDr;
input  [18:0]  BIST_c405dcuBistModeRegIn;
output [18:0]  C405_bistdcuBistModeRegOut;

input          BIST_c405icuBistMbRun;

input  [3:0]   BIST_c405icuBistDebugSi;
input  [3:0]   BIST_c405icuBistDebugEn;
output [3:0]   C405_bisticuBistDebugSo;

input          BIST_c405icuBistShiftDr;
input          BIST_c405icuBistModeRegSi;
output         C405_bisticuBistModeRegSo;

input          BIST_c405icuBistParallelDr;
input  [18:0]  BIST_c405icuBistModeRegIn;
output [18:0]  C405_bisticuBistModeRegOut;


`ifdef VMC_RUN
p405s_vmcmodel PPC405D4 (
`else
PPC405F5V1 PPC405D4(
`endif
     .C405APUDCDHOLD(     C405_apuDcdHold),
     .C405APUDCDFULL(     C405_apuDcdFull),
     .C405APUDCDINSTRUCTION00(     C405_apuDcdInstruction[0]),
     .C405APUDCDINSTRUCTION01(     C405_apuDcdInstruction[1]),
     .C405APUDCDINSTRUCTION02(     C405_apuDcdInstruction[2]),
     .C405APUDCDINSTRUCTION03(     C405_apuDcdInstruction[3]),
     .C405APUDCDINSTRUCTION04(     C405_apuDcdInstruction[4]),
     .C405APUDCDINSTRUCTION05(     C405_apuDcdInstruction[5]),
     .C405APUDCDINSTRUCTION06(     C405_apuDcdInstruction[6]),
     .C405APUDCDINSTRUCTION07(     C405_apuDcdInstruction[7]),
     .C405APUDCDINSTRUCTION08(     C405_apuDcdInstruction[8]),
     .C405APUDCDINSTRUCTION09(     C405_apuDcdInstruction[9]),
     .C405APUDCDINSTRUCTION10(     C405_apuDcdInstruction[10]),
     .C405APUDCDINSTRUCTION11(     C405_apuDcdInstruction[11]),
     .C405APUDCDINSTRUCTION12(     C405_apuDcdInstruction[12]),
     .C405APUDCDINSTRUCTION13(     C405_apuDcdInstruction[13]),
     .C405APUDCDINSTRUCTION14(     C405_apuDcdInstruction[14]),
     .C405APUDCDINSTRUCTION15(     C405_apuDcdInstruction[15]),
     .C405APUDCDINSTRUCTION16(     C405_apuDcdInstruction[16]),
     .C405APUDCDINSTRUCTION17(     C405_apuDcdInstruction[17]),
     .C405APUDCDINSTRUCTION18(     C405_apuDcdInstruction[18]),
     .C405APUDCDINSTRUCTION19(     C405_apuDcdInstruction[19]),
     .C405APUDCDINSTRUCTION20(     C405_apuDcdInstruction[20]),
     .C405APUDCDINSTRUCTION21(     C405_apuDcdInstruction[21]),
     .C405APUDCDINSTRUCTION22(     C405_apuDcdInstruction[22]),
     .C405APUDCDINSTRUCTION23(     C405_apuDcdInstruction[23]),
     .C405APUDCDINSTRUCTION24(     C405_apuDcdInstruction[24]),
     .C405APUDCDINSTRUCTION25(     C405_apuDcdInstruction[25]),
     .C405APUDCDINSTRUCTION26(     C405_apuDcdInstruction[26]),
     .C405APUDCDINSTRUCTION27(     C405_apuDcdInstruction[27]),
     .C405APUDCDINSTRUCTION28(     C405_apuDcdInstruction[28]),
     .C405APUDCDINSTRUCTION29(     C405_apuDcdInstruction[29]),
     .C405APUDCDINSTRUCTION30(     C405_apuDcdInstruction[30]),
     .C405APUDCDINSTRUCTION31(     C405_apuDcdInstruction[31]),
     .C405APUEXEFLUSH(             C405_apuExeFlush),
     .C405APUEXEHOLD(              C405_apuExeHold),
     .C405APUEXELOADDBUS00(        C405_apuExeLoadDBus[0]),
     .C405APUEXELOADDBUS01(        C405_apuExeLoadDBus[1]),
     .C405APUEXELOADDBUS02(        C405_apuExeLoadDBus[2]),
     .C405APUEXELOADDBUS03(        C405_apuExeLoadDBus[3]),
     .C405APUEXELOADDBUS04(        C405_apuExeLoadDBus[4]),
     .C405APUEXELOADDBUS05(        C405_apuExeLoadDBus[5]),
     .C405APUEXELOADDBUS06(        C405_apuExeLoadDBus[6]),
     .C405APUEXELOADDBUS07(        C405_apuExeLoadDBus[7]),
     .C405APUEXELOADDBUS08(        C405_apuExeLoadDBus[8]),
     .C405APUEXELOADDBUS09(        C405_apuExeLoadDBus[9]),
     .C405APUEXELOADDBUS10(        C405_apuExeLoadDBus[10]),
     .C405APUEXELOADDBUS11(        C405_apuExeLoadDBus[11]),
     .C405APUEXELOADDBUS12(        C405_apuExeLoadDBus[12]),
     .C405APUEXELOADDBUS13(        C405_apuExeLoadDBus[13]),
     .C405APUEXELOADDBUS14(        C405_apuExeLoadDBus[14]),
     .C405APUEXELOADDBUS15(        C405_apuExeLoadDBus[15]),
     .C405APUEXELOADDBUS16(        C405_apuExeLoadDBus[16]),
     .C405APUEXELOADDBUS17(        C405_apuExeLoadDBus[17]),
     .C405APUEXELOADDBUS18(        C405_apuExeLoadDBus[18]),
     .C405APUEXELOADDBUS19(        C405_apuExeLoadDBus[19]),
     .C405APUEXELOADDBUS20(        C405_apuExeLoadDBus[20]),
     .C405APUEXELOADDBUS21(        C405_apuExeLoadDBus[21]),
     .C405APUEXELOADDBUS22(        C405_apuExeLoadDBus[22]),
     .C405APUEXELOADDBUS23(        C405_apuExeLoadDBus[23]),
     .C405APUEXELOADDBUS24(        C405_apuExeLoadDBus[24]),
     .C405APUEXELOADDBUS25(        C405_apuExeLoadDBus[25]),
     .C405APUEXELOADDBUS26(        C405_apuExeLoadDBus[26]),
     .C405APUEXELOADDBUS27(        C405_apuExeLoadDBus[27]),
     .C405APUEXELOADDBUS28(        C405_apuExeLoadDBus[28]),
     .C405APUEXELOADDBUS29(        C405_apuExeLoadDBus[29]),
     .C405APUEXELOADDBUS30(        C405_apuExeLoadDBus[30]),
     .C405APUEXELOADDBUS31(        C405_apuExeLoadDBus[31]),
     .C405APUEXELOADDVALID(        C405_apuExeLoadDValid),
     .C405APUEXERADATA00(          C405_apuExeRaData[0]),
     .C405APUEXERADATA01(          C405_apuExeRaData[1]),
     .C405APUEXERADATA02(          C405_apuExeRaData[2]),
     .C405APUEXERADATA03(          C405_apuExeRaData[3]),
     .C405APUEXERADATA04(          C405_apuExeRaData[4]),
     .C405APUEXERADATA05(          C405_apuExeRaData[5]),
     .C405APUEXERADATA06(          C405_apuExeRaData[6]),
     .C405APUEXERADATA07(          C405_apuExeRaData[7]),
     .C405APUEXERADATA08(          C405_apuExeRaData[8]),
     .C405APUEXERADATA09(          C405_apuExeRaData[9]),
     .C405APUEXERADATA10(          C405_apuExeRaData[10]),
     .C405APUEXERADATA11(          C405_apuExeRaData[11]),
     .C405APUEXERADATA12(          C405_apuExeRaData[12]),
     .C405APUEXERADATA13(          C405_apuExeRaData[13]),
     .C405APUEXERADATA14(          C405_apuExeRaData[14]),
     .C405APUEXERADATA15(          C405_apuExeRaData[15]),
     .C405APUEXERADATA16(          C405_apuExeRaData[16]),
     .C405APUEXERADATA17(          C405_apuExeRaData[17]),
     .C405APUEXERADATA18(          C405_apuExeRaData[18]),
     .C405APUEXERADATA19(          C405_apuExeRaData[19]),
     .C405APUEXERADATA20(          C405_apuExeRaData[20]),
     .C405APUEXERADATA21(          C405_apuExeRaData[21]),
     .C405APUEXERADATA22(          C405_apuExeRaData[22]),
     .C405APUEXERADATA23(          C405_apuExeRaData[23]),
     .C405APUEXERADATA24(          C405_apuExeRaData[24]),
     .C405APUEXERADATA25(          C405_apuExeRaData[25]),
     .C405APUEXERADATA26(          C405_apuExeRaData[26]),
     .C405APUEXERADATA27(          C405_apuExeRaData[27]),
     .C405APUEXERADATA28(          C405_apuExeRaData[28]),
     .C405APUEXERADATA29(          C405_apuExeRaData[29]),
     .C405APUEXERADATA30(          C405_apuExeRaData[30]),
     .C405APUEXERADATA31(          C405_apuExeRaData[31]),
     .C405APUEXERBDATA00(          C405_apuExeRbData[0]),
     .C405APUEXERBDATA01(          C405_apuExeRbData[1]),
     .C405APUEXERBDATA02(          C405_apuExeRbData[2]),
     .C405APUEXERBDATA03(          C405_apuExeRbData[3]),
     .C405APUEXERBDATA04(          C405_apuExeRbData[4]),
     .C405APUEXERBDATA05(          C405_apuExeRbData[5]),
     .C405APUEXERBDATA06(          C405_apuExeRbData[6]),
     .C405APUEXERBDATA07(          C405_apuExeRbData[7]),
     .C405APUEXERBDATA08(          C405_apuExeRbData[8]),
     .C405APUEXERBDATA09(          C405_apuExeRbData[9]),
     .C405APUEXERBDATA10(          C405_apuExeRbData[10]),
     .C405APUEXERBDATA11(          C405_apuExeRbData[11]),
     .C405APUEXERBDATA12(          C405_apuExeRbData[12]),
     .C405APUEXERBDATA13(          C405_apuExeRbData[13]),
     .C405APUEXERBDATA14(          C405_apuExeRbData[14]),
     .C405APUEXERBDATA15(          C405_apuExeRbData[15]),
     .C405APUEXERBDATA16(          C405_apuExeRbData[16]),
     .C405APUEXERBDATA17(          C405_apuExeRbData[17]),
     .C405APUEXERBDATA18(          C405_apuExeRbData[18]),
     .C405APUEXERBDATA19(          C405_apuExeRbData[19]),
     .C405APUEXERBDATA20(          C405_apuExeRbData[20]),
     .C405APUEXERBDATA21(          C405_apuExeRbData[21]),
     .C405APUEXERBDATA22(          C405_apuExeRbData[22]),
     .C405APUEXERBDATA23(          C405_apuExeRbData[23]),
     .C405APUEXERBDATA24(          C405_apuExeRbData[24]),
     .C405APUEXERBDATA25(          C405_apuExeRbData[25]),
     .C405APUEXERBDATA26(          C405_apuExeRbData[26]),
     .C405APUEXERBDATA27(          C405_apuExeRbData[27]),
     .C405APUEXERBDATA28(          C405_apuExeRbData[28]),
     .C405APUEXERBDATA29(          C405_apuExeRbData[29]),
     .C405APUEXERBDATA30(          C405_apuExeRbData[30]),
     .C405APUEXERBDATA31(          C405_apuExeRbData[31]),
     .C405APUEXEWDCNT0(            C405_apuExeWdCnt[0]),
     .C405APUEXEWDCNT1(            C405_apuExeWdCnt[1]),
     .C405APUMSRFE0(               C405_apuMsrFE0),
     .C405APUMSRFE1(               C405_apuMsrFE1),
     .C405APUWBBYTEEN0(            C405_apuWbByteEn[0]),
     .C405APUWBBYTEEN1(            C405_apuWbByteEn[1]),
     .C405APUWBBYTEEN2(            C405_apuWbByteEn[2]),
     .C405APUWBBYTEEN3(            C405_apuWbByteEn[3]),
     .C405APUWBENDIAN(             C405_apuWbEndian),
     .C405APUWBFLUSH(              C405_apuWbFlush),
     .C405APUWBHOLD(               C405_apuWbHold),
     .C405APUXERCA(                C405_apuXerCA),
     .C405CPMCORESLEEPREQ(         C405_cpmCoreSleepReq),
     .C405CPMMSRCE(                C405_cpmMsrCE),
     .C405CPMMSREE(                C405_cpmMsrEE),
     .C405CPMTIMERIRQ(             C405_cpmTimerIRQ),
     .C405CPMTIMERRESETREQ(        C405_cpmTimerResetReq),
     .C405DBGLOADDATAONAPUDBUS(    C405_dbgLoadDataOnApuDBus),
     .C405DBGMSRWE(                C405_dbgMsrWE),
     .C405DBGSTOPACK(              C405_dbgStopAck),
     .C405DBGWBCOMPLETE(           C405_dbgWbComplete),
     .C405DBGWBFULL(               C405_dbgWbFull),
     .C405DBGWBIAR00(              C405_dbgWbIar[0]),
     .C405DBGWBIAR01(              C405_dbgWbIar[1]),
     .C405DBGWBIAR02(              C405_dbgWbIar[2]),
     .C405DBGWBIAR03(              C405_dbgWbIar[3]),
     .C405DBGWBIAR04(              C405_dbgWbIar[4]),
     .C405DBGWBIAR05(              C405_dbgWbIar[5]),
     .C405DBGWBIAR06(              C405_dbgWbIar[6]),
     .C405DBGWBIAR07(              C405_dbgWbIar[7]),
     .C405DBGWBIAR08(              C405_dbgWbIar[8]),
     .C405DBGWBIAR09(              C405_dbgWbIar[9]),
     .C405DBGWBIAR10(              C405_dbgWbIar[10]),
     .C405DBGWBIAR11(              C405_dbgWbIar[11]),
     .C405DBGWBIAR12(              C405_dbgWbIar[12]),
     .C405DBGWBIAR13(              C405_dbgWbIar[13]),
     .C405DBGWBIAR14(              C405_dbgWbIar[14]),
     .C405DBGWBIAR15(              C405_dbgWbIar[15]),
     .C405DBGWBIAR16(              C405_dbgWbIar[16]),
     .C405DBGWBIAR17(              C405_dbgWbIar[17]),
     .C405DBGWBIAR18(              C405_dbgWbIar[18]),
     .C405DBGWBIAR19(              C405_dbgWbIar[19]),
     .C405DBGWBIAR20(              C405_dbgWbIar[20]),
     .C405DBGWBIAR21(              C405_dbgWbIar[21]),
     .C405DBGWBIAR22(              C405_dbgWbIar[22]),
     .C405DBGWBIAR23(              C405_dbgWbIar[23]),
     .C405DBGWBIAR24(              C405_dbgWbIar[24]),
     .C405DBGWBIAR25(              C405_dbgWbIar[25]),
     .C405DBGWBIAR26(              C405_dbgWbIar[26]),
     .C405DBGWBIAR27(              C405_dbgWbIar[27]),
     .C405DBGWBIAR28(              C405_dbgWbIar[28]),
     .C405DBGWBIAR29(              C405_dbgWbIar[29]),
     .C405DCRABUS0(                C405_dcrABus[0]),
     .C405DCRABUS1(                C405_dcrABus[1]),
     .C405DCRABUS2(                C405_dcrABus[2]),
     .C405DCRABUS3(                C405_dcrABus[3]),
     .C405DCRABUS4(                C405_dcrABus[4]),
     .C405DCRABUS5(                C405_dcrABus[5]),
     .C405DCRABUS6(                C405_dcrABus[6]),
     .C405DCRABUS7(                C405_dcrABus[7]),
     .C405DCRABUS8(                C405_dcrABus[8]),
     .C405DCRABUS9(                C405_dcrABus[9]),
     .C405DCRDBUSOUT00(            C405_dcrDBusOut[0]),
     .C405DCRDBUSOUT01(            C405_dcrDBusOut[1]),
     .C405DCRDBUSOUT02(            C405_dcrDBusOut[2]),
     .C405DCRDBUSOUT03(            C405_dcrDBusOut[3]),
     .C405DCRDBUSOUT04(            C405_dcrDBusOut[4]),
     .C405DCRDBUSOUT05(            C405_dcrDBusOut[5]),
     .C405DCRDBUSOUT06(            C405_dcrDBusOut[6]),
     .C405DCRDBUSOUT07(            C405_dcrDBusOut[7]),
     .C405DCRDBUSOUT08(            C405_dcrDBusOut[8]),
     .C405DCRDBUSOUT09(            C405_dcrDBusOut[9]),
     .C405DCRDBUSOUT10(            C405_dcrDBusOut[10]),
     .C405DCRDBUSOUT11(            C405_dcrDBusOut[11]),
     .C405DCRDBUSOUT12(            C405_dcrDBusOut[12]),
     .C405DCRDBUSOUT13(            C405_dcrDBusOut[13]),
     .C405DCRDBUSOUT14(            C405_dcrDBusOut[14]),
     .C405DCRDBUSOUT15(            C405_dcrDBusOut[15]),
     .C405DCRDBUSOUT16(            C405_dcrDBusOut[16]),
     .C405DCRDBUSOUT17(            C405_dcrDBusOut[17]),
     .C405DCRDBUSOUT18(            C405_dcrDBusOut[18]),
     .C405DCRDBUSOUT19(            C405_dcrDBusOut[19]),
     .C405DCRDBUSOUT20(            C405_dcrDBusOut[20]),
     .C405DCRDBUSOUT21(            C405_dcrDBusOut[21]),
     .C405DCRDBUSOUT22(            C405_dcrDBusOut[22]),
     .C405DCRDBUSOUT23(            C405_dcrDBusOut[23]),
     .C405DCRDBUSOUT24(            C405_dcrDBusOut[24]),
     .C405DCRDBUSOUT25(            C405_dcrDBusOut[25]),
     .C405DCRDBUSOUT26(            C405_dcrDBusOut[26]),
     .C405DCRDBUSOUT27(            C405_dcrDBusOut[27]),
     .C405DCRDBUSOUT28(            C405_dcrDBusOut[28]),
     .C405DCRDBUSOUT29(            C405_dcrDBusOut[29]),
     .C405DCRDBUSOUT30(            C405_dcrDBusOut[30]),
     .C405DCRDBUSOUT31(            C405_dcrDBusOut[31]),
     .C405DCRREAD(                 C405_dcrRead),
     .C405DCRWRITE(                C405_dcrWrite),
     .C405DSOCMABORTOP(            C405_dsocmAbortOp),
     .C405DSOCMABORTREQ(           C405_dsocmAbortReq),
     .C405DSOCMABUS00(             C405_dsocmABus[0]),
     .C405DSOCMABUS01(             C405_dsocmABus[1]),
     .C405DSOCMABUS02(             C405_dsocmABus[2]),
     .C405DSOCMABUS03(             C405_dsocmABus[3]),
     .C405DSOCMABUS04(             C405_dsocmABus[4]),
     .C405DSOCMABUS05(             C405_dsocmABus[5]),
     .C405DSOCMABUS06(             C405_dsocmABus[6]),
     .C405DSOCMABUS07(             C405_dsocmABus[7]),
     .C405DSOCMABUS08(             C405_dsocmABus[8]),
     .C405DSOCMABUS09(             C405_dsocmABus[9]),
     .C405DSOCMABUS10(             C405_dsocmABus[10]),
     .C405DSOCMABUS11(             C405_dsocmABus[11]),
     .C405DSOCMABUS12(             C405_dsocmABus[12]),
     .C405DSOCMABUS13(             C405_dsocmABus[13]),
     .C405DSOCMABUS14(             C405_dsocmABus[14]),
     .C405DSOCMABUS15(             C405_dsocmABus[15]),
     .C405DSOCMABUS16(             C405_dsocmABus[16]),
     .C405DSOCMABUS17(             C405_dsocmABus[17]),
     .C405DSOCMABUS18(             C405_dsocmABus[18]),
     .C405DSOCMABUS19(             C405_dsocmABus[19]),
     .C405DSOCMABUS20(             C405_dsocmABus[20]),
     .C405DSOCMABUS21(             C405_dsocmABus[21]),
     .C405DSOCMABUS22(             C405_dsocmABus[22]),
     .C405DSOCMABUS23(             C405_dsocmABus[23]),
     .C405DSOCMABUS24(             C405_dsocmABus[24]),
     .C405DSOCMABUS25(             C405_dsocmABus[25]),
     .C405DSOCMABUS26(             C405_dsocmABus[26]),
     .C405DSOCMABUS27(             C405_dsocmABus[27]),
     .C405DSOCMABUS28(             C405_dsocmABus[28]),
     .C405DSOCMABUS29(             C405_dsocmABus[29]),
     .C405DSOCMBYTEEN0(            C405_dsocmByteEn[0]),
     .C405DSOCMBYTEEN1(            C405_dsocmByteEn[1]),
     .C405DSOCMBYTEEN2(            C405_dsocmByteEn[2]),
     .C405DSOCMBYTEEN3(            C405_dsocmByteEn[3]),
     .C405DSOCMCACHEABLE(          C405_dsocmCacheable),
     .C405DSOCMGUARDED(            C405_dsocmGuarded),
     .C405DSOCMLOADREQ(            C405_dsocmLoadReq),
     .C405DSOCMSTOREREQ(           C405_dsocmStoreReq),
     .C405DSOCMSTRINGMULTIPLE(     C405_dsocmStringMultiple),
     .C405DSOCMU0ATTR(             C405_dsocmU0Attr),
     .C405DSOCMWAIT(               C405_dsocmWait),
     .C405DSOCMWRDBUS00(           C405_dsocmWrDBus[0]),
     .C405DSOCMWRDBUS01(           C405_dsocmWrDBus[1]),
     .C405DSOCMWRDBUS02(           C405_dsocmWrDBus[2]),
     .C405DSOCMWRDBUS03(           C405_dsocmWrDBus[3]),
     .C405DSOCMWRDBUS04(           C405_dsocmWrDBus[4]),
     .C405DSOCMWRDBUS05(           C405_dsocmWrDBus[5]),
     .C405DSOCMWRDBUS06(           C405_dsocmWrDBus[6]),
     .C405DSOCMWRDBUS07(           C405_dsocmWrDBus[7]),
     .C405DSOCMWRDBUS08(           C405_dsocmWrDBus[8]),
     .C405DSOCMWRDBUS09(           C405_dsocmWrDBus[9]),
     .C405DSOCMWRDBUS10(           C405_dsocmWrDBus[10]),
     .C405DSOCMWRDBUS11(           C405_dsocmWrDBus[11]),
     .C405DSOCMWRDBUS12(           C405_dsocmWrDBus[12]),
     .C405DSOCMWRDBUS13(           C405_dsocmWrDBus[13]),
     .C405DSOCMWRDBUS14(           C405_dsocmWrDBus[14]),
     .C405DSOCMWRDBUS15(           C405_dsocmWrDBus[15]),
     .C405DSOCMWRDBUS16(           C405_dsocmWrDBus[16]),
     .C405DSOCMWRDBUS17(           C405_dsocmWrDBus[17]),
     .C405DSOCMWRDBUS18(           C405_dsocmWrDBus[18]),
     .C405DSOCMWRDBUS19(           C405_dsocmWrDBus[19]),
     .C405DSOCMWRDBUS20(           C405_dsocmWrDBus[20]),
     .C405DSOCMWRDBUS21(           C405_dsocmWrDBus[21]),
     .C405DSOCMWRDBUS22(           C405_dsocmWrDBus[22]),
     .C405DSOCMWRDBUS23(           C405_dsocmWrDBus[23]),
     .C405DSOCMWRDBUS24(           C405_dsocmWrDBus[24]),
     .C405DSOCMWRDBUS25(           C405_dsocmWrDBus[25]),
     .C405DSOCMWRDBUS26(           C405_dsocmWrDBus[26]),
     .C405DSOCMWRDBUS27(           C405_dsocmWrDBus[27]),
     .C405DSOCMWRDBUS28(           C405_dsocmWrDBus[28]),
     .C405DSOCMWRDBUS29(           C405_dsocmWrDBus[29]),
     .C405DSOCMWRDBUS30(           C405_dsocmWrDBus[30]),
     .C405DSOCMWRDBUS31(           C405_dsocmWrDBus[31]),
     .C405DSOCMXLATEVALID(         C405_dsocmXlateValid),
     .C405ISOCMABORT(              C405_isocmAbort),
     .C405ISOCMABUS00(             C405_isocmABus[0]),
     .C405ISOCMABUS01(             C405_isocmABus[1]),
     .C405ISOCMABUS02(             C405_isocmABus[2]),
     .C405ISOCMABUS03(             C405_isocmABus[3]),
     .C405ISOCMABUS04(             C405_isocmABus[4]),
     .C405ISOCMABUS05(             C405_isocmABus[5]),
     .C405ISOCMABUS06(             C405_isocmABus[6]),
     .C405ISOCMABUS07(             C405_isocmABus[7]),
     .C405ISOCMABUS08(             C405_isocmABus[8]),
     .C405ISOCMABUS09(             C405_isocmABus[9]),
     .C405ISOCMABUS10(             C405_isocmABus[10]),
     .C405ISOCMABUS11(             C405_isocmABus[11]),
     .C405ISOCMABUS12(             C405_isocmABus[12]),
     .C405ISOCMABUS13(             C405_isocmABus[13]),
     .C405ISOCMABUS14(             C405_isocmABus[14]),
     .C405ISOCMABUS15(             C405_isocmABus[15]),
     .C405ISOCMABUS16(             C405_isocmABus[16]),
     .C405ISOCMABUS17(             C405_isocmABus[17]),
     .C405ISOCMABUS18(             C405_isocmABus[18]),
     .C405ISOCMABUS19(             C405_isocmABus[19]),
     .C405ISOCMABUS20(             C405_isocmABus[20]),
     .C405ISOCMABUS21(             C405_isocmABus[21]),
     .C405ISOCMABUS22(             C405_isocmABus[22]),
     .C405ISOCMABUS23(             C405_isocmABus[23]),
     .C405ISOCMABUS24(             C405_isocmABus[24]),
     .C405ISOCMABUS25(             C405_isocmABus[25]),
     .C405ISOCMABUS26(             C405_isocmABus[26]),
     .C405ISOCMABUS27(             C405_isocmABus[27]),
     .C405ISOCMABUS28(             C405_isocmABus[28]),
     .C405ISOCMABUS29(             C405_isocmABus[29]),
     .C405ISOCMCACHEABLE(          C405_isocmCacheable),
     .C405ISOCMCONTEXTSYNC(        C405_isocmContextSync),
     .C405ISOCMICUREADY(           C405_isocmIcuReady),
     .C405ISOCMREQPENDING(         C405_isocmReqPending),
     .C405ISOCMU0ATTR(             C405_isocmU0Attr),
     .C405ISOCMXLATEVALID(         C405_isocmXlateValid),
     .C405JTGCAPTUREDR(            C405_jtgCaptureDR),
     .C405JTGEXTEST(               C405_jtgExtest),
     .C405JTGPGMOUT(               C405_jtgPgmOut),
     .C405JTGSHIFTDR(              C405_jtgShiftDR),
     .C405JTGTDO(                  C405_jtgTDO),
     .C405JTGTDOEN(                C405_jtgTDOEn),
     .C405JTGUPDATEDR(             C405_jtgUpdateDR),
     .C405TESTDIAGABISTDONE(       C405_testDiagAbistDone),
     .C405PLBDCUABORT(             C405_plbDcuAbort),
     .C405PLBDCUABUS00(            C405_plbDcuABus[0]),
     .C405PLBDCUABUS01(            C405_plbDcuABus[1]),
     .C405PLBDCUABUS02(            C405_plbDcuABus[2]),
     .C405PLBDCUABUS03(            C405_plbDcuABus[3]),
     .C405PLBDCUABUS04(            C405_plbDcuABus[4]),
     .C405PLBDCUABUS05(            C405_plbDcuABus[5]),
     .C405PLBDCUABUS06(            C405_plbDcuABus[6]),
     .C405PLBDCUABUS07(            C405_plbDcuABus[7]),
     .C405PLBDCUABUS08(            C405_plbDcuABus[8]),
     .C405PLBDCUABUS09(            C405_plbDcuABus[9]),
     .C405PLBDCUABUS10(            C405_plbDcuABus[10]),
     .C405PLBDCUABUS11(            C405_plbDcuABus[11]),
     .C405PLBDCUABUS12(            C405_plbDcuABus[12]),
     .C405PLBDCUABUS13(            C405_plbDcuABus[13]),
     .C405PLBDCUABUS14(            C405_plbDcuABus[14]),
     .C405PLBDCUABUS15(            C405_plbDcuABus[15]),
     .C405PLBDCUABUS16(            C405_plbDcuABus[16]),
     .C405PLBDCUABUS17(            C405_plbDcuABus[17]),
     .C405PLBDCUABUS18(            C405_plbDcuABus[18]),
     .C405PLBDCUABUS19(            C405_plbDcuABus[19]),
     .C405PLBDCUABUS20(            C405_plbDcuABus[20]),
     .C405PLBDCUABUS21(            C405_plbDcuABus[21]),
     .C405PLBDCUABUS22(            C405_plbDcuABus[22]),
     .C405PLBDCUABUS23(            C405_plbDcuABus[23]),
     .C405PLBDCUABUS24(            C405_plbDcuABus[24]),
     .C405PLBDCUABUS25(            C405_plbDcuABus[25]),
     .C405PLBDCUABUS26(            C405_plbDcuABus[26]),
     .C405PLBDCUABUS27(            C405_plbDcuABus[27]),
     .C405PLBDCUABUS28(            C405_plbDcuABus[28]),
     .C405PLBDCUABUS29(            C405_plbDcuABus[29]),
     .C405PLBDCUABUS30(            C405_plbDcuABus[30]),
     .C405PLBDCUABUS31(            C405_plbDcuABus[31]),
     .C405PLBDCUBE0(               C405_plbDcuBE[0]),
     .C405PLBDCUBE1(               C405_plbDcuBE[1]),
     .C405PLBDCUBE2(               C405_plbDcuBE[2]),
     .C405PLBDCUBE3(               C405_plbDcuBE[3]),
     .C405PLBDCUBE4(               C405_plbDcuBE[4]),
     .C405PLBDCUBE5(               C405_plbDcuBE[5]),
     .C405PLBDCUBE6(               C405_plbDcuBE[6]),
     .C405PLBDCUBE7(               C405_plbDcuBE[7]),
     .C405PLBDCUCACHEABLE(         C405_plbDcuCacheable),
     .C405PLBDCUGUARDED(           C405_plbDcuGuarded),
     .C405PLBDCUPRIORITY0(         C405_plbDcuPriority[0]),
     .C405PLBDCUPRIORITY1(         C405_plbDcuPriority[1]),
     .C405PLBDCUREQUEST(           C405_plbDcuRequest),
     .C405PLBDCURNW(               C405_plbDcuRNW),
     .C405PLBDCUSIZE2(             C405_plbDcuSize2),
     .C405PLBDCUU0ATTR(            C405_plbDcuU0Attr),
     .C405PLBDCUWRDBUS00(          C405_plbDcuWrDBus[0]),
     .C405PLBDCUWRDBUS01(          C405_plbDcuWrDBus[1]),
     .C405PLBDCUWRDBUS02(          C405_plbDcuWrDBus[2]),
     .C405PLBDCUWRDBUS03(          C405_plbDcuWrDBus[3]),
     .C405PLBDCUWRDBUS04(          C405_plbDcuWrDBus[4]),
     .C405PLBDCUWRDBUS05(          C405_plbDcuWrDBus[5]),
     .C405PLBDCUWRDBUS06(          C405_plbDcuWrDBus[6]),
     .C405PLBDCUWRDBUS07(          C405_plbDcuWrDBus[7]),
     .C405PLBDCUWRDBUS08(          C405_plbDcuWrDBus[8]),
     .C405PLBDCUWRDBUS09(          C405_plbDcuWrDBus[9]),
     .C405PLBDCUWRDBUS10(          C405_plbDcuWrDBus[10]),
     .C405PLBDCUWRDBUS11(          C405_plbDcuWrDBus[11]),
     .C405PLBDCUWRDBUS12(          C405_plbDcuWrDBus[12]),
     .C405PLBDCUWRDBUS13(          C405_plbDcuWrDBus[13]),
     .C405PLBDCUWRDBUS14(          C405_plbDcuWrDBus[14]),
     .C405PLBDCUWRDBUS15(          C405_plbDcuWrDBus[15]),
     .C405PLBDCUWRDBUS16(          C405_plbDcuWrDBus[16]),
     .C405PLBDCUWRDBUS17(          C405_plbDcuWrDBus[17]),
     .C405PLBDCUWRDBUS18(          C405_plbDcuWrDBus[18]),
     .C405PLBDCUWRDBUS19(          C405_plbDcuWrDBus[19]),
     .C405PLBDCUWRDBUS20(          C405_plbDcuWrDBus[20]),
     .C405PLBDCUWRDBUS21(          C405_plbDcuWrDBus[21]),
     .C405PLBDCUWRDBUS22(          C405_plbDcuWrDBus[22]),
     .C405PLBDCUWRDBUS23(          C405_plbDcuWrDBus[23]),
     .C405PLBDCUWRDBUS24(          C405_plbDcuWrDBus[24]),
     .C405PLBDCUWRDBUS25(          C405_plbDcuWrDBus[25]),
     .C405PLBDCUWRDBUS26(          C405_plbDcuWrDBus[26]),
     .C405PLBDCUWRDBUS27(          C405_plbDcuWrDBus[27]),
     .C405PLBDCUWRDBUS28(          C405_plbDcuWrDBus[28]),
     .C405PLBDCUWRDBUS29(          C405_plbDcuWrDBus[29]),
     .C405PLBDCUWRDBUS30(          C405_plbDcuWrDBus[30]),
     .C405PLBDCUWRDBUS31(          C405_plbDcuWrDBus[31]),
     .C405PLBDCUWRDBUS32(          C405_plbDcuWrDBus[32]),
     .C405PLBDCUWRDBUS33(          C405_plbDcuWrDBus[33]),
     .C405PLBDCUWRDBUS34(          C405_plbDcuWrDBus[34]),
     .C405PLBDCUWRDBUS35(          C405_plbDcuWrDBus[35]),
     .C405PLBDCUWRDBUS36(          C405_plbDcuWrDBus[36]),
     .C405PLBDCUWRDBUS37(          C405_plbDcuWrDBus[37]),
     .C405PLBDCUWRDBUS38(          C405_plbDcuWrDBus[38]),
     .C405PLBDCUWRDBUS39(          C405_plbDcuWrDBus[39]),
     .C405PLBDCUWRDBUS40(          C405_plbDcuWrDBus[40]),
     .C405PLBDCUWRDBUS41(          C405_plbDcuWrDBus[41]),
     .C405PLBDCUWRDBUS42(          C405_plbDcuWrDBus[42]),
     .C405PLBDCUWRDBUS43(          C405_plbDcuWrDBus[43]),
     .C405PLBDCUWRDBUS44(          C405_plbDcuWrDBus[44]),
     .C405PLBDCUWRDBUS45(          C405_plbDcuWrDBus[45]),
     .C405PLBDCUWRDBUS46(          C405_plbDcuWrDBus[46]),
     .C405PLBDCUWRDBUS47(          C405_plbDcuWrDBus[47]),
     .C405PLBDCUWRDBUS48(          C405_plbDcuWrDBus[48]),
     .C405PLBDCUWRDBUS49(          C405_plbDcuWrDBus[49]),
     .C405PLBDCUWRDBUS50(          C405_plbDcuWrDBus[50]),
     .C405PLBDCUWRDBUS51(          C405_plbDcuWrDBus[51]),
     .C405PLBDCUWRDBUS52(          C405_plbDcuWrDBus[52]),
     .C405PLBDCUWRDBUS53(          C405_plbDcuWrDBus[53]),
     .C405PLBDCUWRDBUS54(          C405_plbDcuWrDBus[54]),
     .C405PLBDCUWRDBUS55(          C405_plbDcuWrDBus[55]),
     .C405PLBDCUWRDBUS56(          C405_plbDcuWrDBus[56]),
     .C405PLBDCUWRDBUS57(          C405_plbDcuWrDBus[57]),
     .C405PLBDCUWRDBUS58(          C405_plbDcuWrDBus[58]),
     .C405PLBDCUWRDBUS59(          C405_plbDcuWrDBus[59]),
     .C405PLBDCUWRDBUS60(          C405_plbDcuWrDBus[60]),
     .C405PLBDCUWRDBUS61(          C405_plbDcuWrDBus[61]),
     .C405PLBDCUWRDBUS62(          C405_plbDcuWrDBus[62]),
     .C405PLBDCUWRDBUS63(          C405_plbDcuWrDBus[63]),
     .C405PLBDCUWRITETHRU(         C405_plbDcuWriteThru),
     .C405PLBICUABORT(             C405_plbIcuAbort),
     .C405PLBICUABUS00(            C405_plbIcuABus[0]),
     .C405PLBICUABUS01(            C405_plbIcuABus[1]),
     .C405PLBICUABUS02(            C405_plbIcuABus[2]),
     .C405PLBICUABUS03(            C405_plbIcuABus[3]),
     .C405PLBICUABUS04(            C405_plbIcuABus[4]),
     .C405PLBICUABUS05(            C405_plbIcuABus[5]),
     .C405PLBICUABUS06(            C405_plbIcuABus[6]),
     .C405PLBICUABUS07(            C405_plbIcuABus[7]),
     .C405PLBICUABUS08(            C405_plbIcuABus[8]),
     .C405PLBICUABUS09(            C405_plbIcuABus[9]),
     .C405PLBICUABUS10(            C405_plbIcuABus[10]),
     .C405PLBICUABUS11(            C405_plbIcuABus[11]),
     .C405PLBICUABUS12(            C405_plbIcuABus[12]),
     .C405PLBICUABUS13(            C405_plbIcuABus[13]),
     .C405PLBICUABUS14(            C405_plbIcuABus[14]),
     .C405PLBICUABUS15(            C405_plbIcuABus[15]),
     .C405PLBICUABUS16(            C405_plbIcuABus[16]),
     .C405PLBICUABUS17(            C405_plbIcuABus[17]),
     .C405PLBICUABUS18(            C405_plbIcuABus[18]),
     .C405PLBICUABUS19(            C405_plbIcuABus[19]),
     .C405PLBICUABUS20(            C405_plbIcuABus[20]),
     .C405PLBICUABUS21(            C405_plbIcuABus[21]),
     .C405PLBICUABUS22(            C405_plbIcuABus[22]),
     .C405PLBICUABUS23(            C405_plbIcuABus[23]),
     .C405PLBICUABUS24(            C405_plbIcuABus[24]),
     .C405PLBICUABUS25(            C405_plbIcuABus[25]),
     .C405PLBICUABUS26(            C405_plbIcuABus[26]),
     .C405PLBICUABUS27(            C405_plbIcuABus[27]),
     .C405PLBICUABUS28(            C405_plbIcuABus[28]),
     .C405PLBICUABUS29(            C405_plbIcuABus[29]),
     .C405PLBICUCACHEABLE(         C405_plbIcuCacheable),
     .C405PLBICUPRIORITY0(         C405_plbIcuPriority[0]),
     .C405PLBICUPRIORITY1(         C405_plbIcuPriority[1]),
     .C405PLBICUREQUEST(           C405_plbIcuRequest),
     .C405PLBICUSIZE2(             C405_plbIcuSize[2]),
     .C405PLBICUSIZE3(             C405_plbIcuSize[3]),
     .C405PLBICUU0ATTR(            C405_plbIcuU0Attr),
     .C405RSTCHIPRESETREQ(         C405_rstChipResetReq),
     .C405RSTCORERESETREQ(         C405_rstCoreResetReq),
     .C405RSTSYSTEMRESETREQ(       C405_rstSystemResetReq),
     .C405TRCCYCLE(                C405_trcCycle),
     .C405TRCEVENEXECUTIONSTATUS0( C405_trcEvenExecutionStatus[0]),
     .C405TRCEVENEXECUTIONSTATUS1( C405_trcEvenExecutionStatus[1]),
     .C405TRCODDEXECUTIONSTATUS0(  C405_trcOddExecutionStatus[0]),
     .C405TRCODDEXECUTIONSTATUS1(  C405_trcOddExecutionStatus[1]),
     .C405TRCTRACESTATUS0(         C405_trcTraceStatus[0]),
     .C405TRCTRACESTATUS1(         C405_trcTraceStatus[1]),
     .C405TRCTRACESTATUS2(         C405_trcTraceStatus[2]),
     .C405TRCTRACESTATUS3(         C405_trcTraceStatus[3]),
     .C405TRCTRIGGEREVENTOUT(      C405_trcTriggerEventOut),
     .C405TRCTRIGGEREVENTTYPE0(    C405_trcTriggerEventType[0]),
     .C405TRCTRIGGEREVENTTYPE1(    C405_trcTriggerEventType[1]),
     .C405TRCTRIGGEREVENTTYPE2(    C405_trcTriggerEventType[2]),
     .C405TRCTRIGGEREVENTTYPE3(    C405_trcTriggerEventType[3]),
     .C405TRCTRIGGEREVENTTYPE4(    C405_trcTriggerEventType[4]),
     .C405TRCTRIGGEREVENTTYPE5(    C405_trcTriggerEventType[5]),
     .C405TRCTRIGGEREVENTTYPE6(    C405_trcTriggerEventType[6]),
     .C405TRCTRIGGEREVENTTYPE7(    C405_trcTriggerEventType[7]),
     .C405TRCTRIGGEREVENTTYPE8(    C405_trcTriggerEventType[8]),
     .C405TRCTRIGGEREVENTTYPE9(    C405_trcTriggerEventType[9]),
     .C405TRCTRIGGEREVENTTYPE10(   C405_trcTriggerEventType[10]),
     .C405XXXMACHINECHECK(         C405_xxxMachineCheck),
     .APUC405DCDAPUOP(             APU_c405DcdApuOp),
     .APUC405DCDCREN(              APU_c405DcdCREn),
     .APUC405DCDFORCEALGN(         APU_c405DcdForceAlgn),
     .APUC405DCDFORCEBESTEERING(   APU_c405DcdForceBESteering),
     .APUC405DCDFPUOP(             APU_c405DcdFpuOp),
     .APUC405DCDGPRWRITE(          APU_c405DcdGprWrite),
     .APUC405DCDLDSTBYTE(          APU_c405DcdLdStByte),
     .APUC405DCDLDSTDW(            APU_c405DcdLdStDw),
     .APUC405DCDLDSTHW(            APU_c405DcdLdStHw),
     .APUC405DCDLDSTQW(            APU_c405DcdLdStQw),
     .APUC405DCDLDSTWD(            APU_c405DcdLdStWd),
     .APUC405DCDLOAD(              APU_c405DcdLoad),
     .APUC405DCDPRIVOP(            APU_c405DcdPrivOp),
     .APUC405DCDRAEN(              APU_c405DcdRaEn),
     .APUC405DCDRBEN(              APU_c405DcdRbEn),
     .APUC405DCDSTORE(             APU_c405DcdStore),
     .APUC405DCDTRAPBE(            APU_c405DcdTrapBE),
     .APUC405DCDTRAPLE(            APU_c405DcdTrapLE),
     .APUC405DCDUPDATE(            APU_c405DcdUpdate),
     .APUC405DCDVALIDOP(           APU_c405DcdValidOp),
     .APUC405DCDXERCAEN(           APU_c405DcdXerCAEn),
     .APUC405DCDXEROVEN(           APU_c405DcdXerOVEn),
     .APUC405EXCEPTION(            APU_c405Exception),
     .APUC405EXEBLOCKINGMCO(       APU_c405ExeBlockingMCO),
     .APUC405EXEBUSY(              APU_c405ExeBusy),
     .APUC405EXECR0(               APU_c405ExeCR[0]),
     .APUC405EXECR1(               APU_c405ExeCR[1]),
     .APUC405EXECR2(               APU_c405ExeCR[2]),
     .APUC405EXECR3(               APU_c405ExeCR[3]),
     .APUC405EXECRFIELD0(          APU_c405ExeCRField[0]),
     .APUC405EXECRFIELD1(          APU_c405ExeCRField[1]),
     .APUC405EXECRFIELD2(          APU_c405ExeCRField[2]),
     .APUC405EXELDDEPEND(          APU_c405ExeLdDepend),
     .APUC405EXENONBLOCKINGMCO(    APU_c405ExeNonBlockingMCO),
     .APUC405EXERESULT00(          APU_c405ExeResult[0]),
     .APUC405EXERESULT01(          APU_c405ExeResult[1]),
     .APUC405EXERESULT02(          APU_c405ExeResult[2]),
     .APUC405EXERESULT03(          APU_c405ExeResult[3]),
     .APUC405EXERESULT04(          APU_c405ExeResult[4]),
     .APUC405EXERESULT05(          APU_c405ExeResult[5]),
     .APUC405EXERESULT06(          APU_c405ExeResult[6]),
     .APUC405EXERESULT07(          APU_c405ExeResult[7]),
     .APUC405EXERESULT08(          APU_c405ExeResult[8]),
     .APUC405EXERESULT09(          APU_c405ExeResult[9]),
     .APUC405EXERESULT10(          APU_c405ExeResult[10]),
     .APUC405EXERESULT11(          APU_c405ExeResult[11]),
     .APUC405EXERESULT12(          APU_c405ExeResult[12]),
     .APUC405EXERESULT13(          APU_c405ExeResult[13]),
     .APUC405EXERESULT14(          APU_c405ExeResult[14]),
     .APUC405EXERESULT15(          APU_c405ExeResult[15]),
     .APUC405EXERESULT16(          APU_c405ExeResult[16]),
     .APUC405EXERESULT17(          APU_c405ExeResult[17]),
     .APUC405EXERESULT18(          APU_c405ExeResult[18]),
     .APUC405EXERESULT19(          APU_c405ExeResult[19]),
     .APUC405EXERESULT20(          APU_c405ExeResult[20]),
     .APUC405EXERESULT21(          APU_c405ExeResult[21]),
     .APUC405EXERESULT22(          APU_c405ExeResult[22]),
     .APUC405EXERESULT23(          APU_c405ExeResult[23]),
     .APUC405EXERESULT24(          APU_c405ExeResult[24]),
     .APUC405EXERESULT25(          APU_c405ExeResult[25]),
     .APUC405EXERESULT26(          APU_c405ExeResult[26]),
     .APUC405EXERESULT27(          APU_c405ExeResult[27]),
     .APUC405EXERESULT28(          APU_c405ExeResult[28]),
     .APUC405EXERESULT29(          APU_c405ExeResult[29]),
     .APUC405EXERESULT30(          APU_c405ExeResult[30]),
     .APUC405EXERESULT31(          APU_c405ExeResult[31]),
     .APUC405EXEXERCA(             APU_c405ExeXerCA),
     .APUC405EXEXEROV(             APU_c405ExeXerOV),
     .APUC405FPUEXCEPTION(         APU_c405FpuException),
     .APUC405LWBLDDEPEND(          APU_c405LwbLdDepend),
     .APUC405SLEEPREQ(             APU_c405SleepReq),
     .APUC405WBLDDEPEND(           APU_c405WbLdDepend),
     .CPMC405CLOCK(                CPM_c405Clock),
     .CPMC405CPUCLKENCCLK(         CPM_c405CpuClkEn_CClk),
     .CPMC405CORECLKINACTIVE(      CPM_c405CoreClkInactive),
     .CPMC405JTAGCLKENCCLK(        CPM_c405JtagClkEn_CClk),
     .CPMC405PLBSAMPLECYCLE(       CPM_c405PlbSampleCycle),
     .CPMC405TIMERCLKENCCLK(       CPM_c405TimerClkEn_CClk),
     .CPMC405TIMERTICK(            CPM_c405TimerTick),
     .DBGC405DEBUGHALT(            DBG_c405DebugHalt),
     .DBGC405EXTBUSHOLDACK(        DBG_c405ExtBusHoldAck),
     .DBGC405UNCONDDEBUGEVENT(     DBG_c405UncondDebugEvent),
     .DCRC405ACK(                  DCR_c405Ack),
     .DCRC405DBUSIN00(             DCR_c405DBusIn[0]),
     .DCRC405DBUSIN01(             DCR_c405DBusIn[1]),
     .DCRC405DBUSIN02(             DCR_c405DBusIn[2]),
     .DCRC405DBUSIN03(             DCR_c405DBusIn[3]),
     .DCRC405DBUSIN04(             DCR_c405DBusIn[4]),
     .DCRC405DBUSIN05(             DCR_c405DBusIn[5]),
     .DCRC405DBUSIN06(             DCR_c405DBusIn[6]),
     .DCRC405DBUSIN07(             DCR_c405DBusIn[7]),
     .DCRC405DBUSIN08(             DCR_c405DBusIn[8]),
     .DCRC405DBUSIN09(             DCR_c405DBusIn[9]),
     .DCRC405DBUSIN10(             DCR_c405DBusIn[10]),
     .DCRC405DBUSIN11(             DCR_c405DBusIn[11]),
     .DCRC405DBUSIN12(             DCR_c405DBusIn[12]),
     .DCRC405DBUSIN13(             DCR_c405DBusIn[13]),
     .DCRC405DBUSIN14(             DCR_c405DBusIn[14]),
     .DCRC405DBUSIN15(             DCR_c405DBusIn[15]),
     .DCRC405DBUSIN16(             DCR_c405DBusIn[16]),
     .DCRC405DBUSIN17(             DCR_c405DBusIn[17]),
     .DCRC405DBUSIN18(             DCR_c405DBusIn[18]),
     .DCRC405DBUSIN19(             DCR_c405DBusIn[19]),
     .DCRC405DBUSIN20(             DCR_c405DBusIn[20]),
     .DCRC405DBUSIN21(             DCR_c405DBusIn[21]),
     .DCRC405DBUSIN22(             DCR_c405DBusIn[22]),
     .DCRC405DBUSIN23(             DCR_c405DBusIn[23]),
     .DCRC405DBUSIN24(             DCR_c405DBusIn[24]),
     .DCRC405DBUSIN25(             DCR_c405DBusIn[25]),
     .DCRC405DBUSIN26(             DCR_c405DBusIn[26]),
     .DCRC405DBUSIN27(             DCR_c405DBusIn[27]),
     .DCRC405DBUSIN28(             DCR_c405DBusIn[28]),
     .DCRC405DBUSIN29(             DCR_c405DBusIn[29]),
     .DCRC405DBUSIN30(             DCR_c405DBusIn[30]),
     .DCRC405DBUSIN31(             DCR_c405DBusIn[31]),
     .DSOCMC405COMPLETE(           DSOCM_c405Complete),
     .DSOCMC405DISOPERANDFWD(      DSOCM_c405DisOperandFwd),
     .DSOCMC405HOLD(               DSOCM_c405Hold),
     .DSOCMC405RDDBUS00(           DSOCM_c405RdDBus[0]),
     .DSOCMC405RDDBUS01(           DSOCM_c405RdDBus[1]),
     .DSOCMC405RDDBUS02(           DSOCM_c405RdDBus[2]),
     .DSOCMC405RDDBUS03(           DSOCM_c405RdDBus[3]),
     .DSOCMC405RDDBUS04(           DSOCM_c405RdDBus[4]),
     .DSOCMC405RDDBUS05(           DSOCM_c405RdDBus[5]),
     .DSOCMC405RDDBUS06(           DSOCM_c405RdDBus[6]),
     .DSOCMC405RDDBUS07(           DSOCM_c405RdDBus[7]),
     .DSOCMC405RDDBUS08(           DSOCM_c405RdDBus[8]),
     .DSOCMC405RDDBUS09(           DSOCM_c405RdDBus[9]),
     .DSOCMC405RDDBUS10(           DSOCM_c405RdDBus[10]),
     .DSOCMC405RDDBUS11(           DSOCM_c405RdDBus[11]),
     .DSOCMC405RDDBUS12(           DSOCM_c405RdDBus[12]),
     .DSOCMC405RDDBUS13(           DSOCM_c405RdDBus[13]),
     .DSOCMC405RDDBUS14(           DSOCM_c405RdDBus[14]),
     .DSOCMC405RDDBUS15(           DSOCM_c405RdDBus[15]),
     .DSOCMC405RDDBUS16(           DSOCM_c405RdDBus[16]),
     .DSOCMC405RDDBUS17(           DSOCM_c405RdDBus[17]),
     .DSOCMC405RDDBUS18(           DSOCM_c405RdDBus[18]),
     .DSOCMC405RDDBUS19(           DSOCM_c405RdDBus[19]),
     .DSOCMC405RDDBUS20(           DSOCM_c405RdDBus[20]),
     .DSOCMC405RDDBUS21(           DSOCM_c405RdDBus[21]),
     .DSOCMC405RDDBUS22(           DSOCM_c405RdDBus[22]),
     .DSOCMC405RDDBUS23(           DSOCM_c405RdDBus[23]),
     .DSOCMC405RDDBUS24(           DSOCM_c405RdDBus[24]),
     .DSOCMC405RDDBUS25(           DSOCM_c405RdDBus[25]),
     .DSOCMC405RDDBUS26(           DSOCM_c405RdDBus[26]),
     .DSOCMC405RDDBUS27(           DSOCM_c405RdDBus[27]),
     .DSOCMC405RDDBUS28(           DSOCM_c405RdDBus[28]),
     .DSOCMC405RDDBUS29(           DSOCM_c405RdDBus[29]),
     .DSOCMC405RDDBUS30(           DSOCM_c405RdDBus[30]),
     .DSOCMC405RDDBUS31(           DSOCM_c405RdDBus[31]),
     .EICC405CRITINPUTIRQ(         EIC_c405CritInputIRQ),
     .EICC405EXTINPUTIRQ(          EIC_c405ExtInputIRQ),
     .ISOCMC405HOLD(               ISOCM_c405Hold),
     .ISOCMC405RDDBUS00(           ISOCM_c405RdDBus[0]),
     .ISOCMC405RDDBUS01(           ISOCM_c405RdDBus[1]),
     .ISOCMC405RDDBUS02(           ISOCM_c405RdDBus[2]),
     .ISOCMC405RDDBUS03(           ISOCM_c405RdDBus[3]),
     .ISOCMC405RDDBUS04(           ISOCM_c405RdDBus[4]),
     .ISOCMC405RDDBUS05(           ISOCM_c405RdDBus[5]),
     .ISOCMC405RDDBUS06(           ISOCM_c405RdDBus[6]),
     .ISOCMC405RDDBUS07(           ISOCM_c405RdDBus[7]),
     .ISOCMC405RDDBUS08(           ISOCM_c405RdDBus[8]),
     .ISOCMC405RDDBUS09(           ISOCM_c405RdDBus[9]),
     .ISOCMC405RDDBUS10(           ISOCM_c405RdDBus[10]),
     .ISOCMC405RDDBUS11(           ISOCM_c405RdDBus[11]),
     .ISOCMC405RDDBUS12(           ISOCM_c405RdDBus[12]),
     .ISOCMC405RDDBUS13(           ISOCM_c405RdDBus[13]),
     .ISOCMC405RDDBUS14(           ISOCM_c405RdDBus[14]),
     .ISOCMC405RDDBUS15(           ISOCM_c405RdDBus[15]),
     .ISOCMC405RDDBUS16(           ISOCM_c405RdDBus[16]),
     .ISOCMC405RDDBUS17(           ISOCM_c405RdDBus[17]),
     .ISOCMC405RDDBUS18(           ISOCM_c405RdDBus[18]),
     .ISOCMC405RDDBUS19(           ISOCM_c405RdDBus[19]),
     .ISOCMC405RDDBUS20(           ISOCM_c405RdDBus[20]),
     .ISOCMC405RDDBUS21(           ISOCM_c405RdDBus[21]),
     .ISOCMC405RDDBUS22(           ISOCM_c405RdDBus[22]),
     .ISOCMC405RDDBUS23(           ISOCM_c405RdDBus[23]),
     .ISOCMC405RDDBUS24(           ISOCM_c405RdDBus[24]),
     .ISOCMC405RDDBUS25(           ISOCM_c405RdDBus[25]),
     .ISOCMC405RDDBUS26(           ISOCM_c405RdDBus[26]),
     .ISOCMC405RDDBUS27(           ISOCM_c405RdDBus[27]),
     .ISOCMC405RDDBUS28(           ISOCM_c405RdDBus[28]),
     .ISOCMC405RDDBUS29(           ISOCM_c405RdDBus[29]),
     .ISOCMC405RDDBUS30(           ISOCM_c405RdDBus[30]),
     .ISOCMC405RDDBUS31(           ISOCM_c405RdDBus[31]),
     .ISOCMC405RDDBUS32(           ISOCM_c405RdDBus[32]),
     .ISOCMC405RDDBUS33(           ISOCM_c405RdDBus[33]),
     .ISOCMC405RDDBUS34(           ISOCM_c405RdDBus[34]),
     .ISOCMC405RDDBUS35(           ISOCM_c405RdDBus[35]),
     .ISOCMC405RDDBUS36(           ISOCM_c405RdDBus[36]),
     .ISOCMC405RDDBUS37(           ISOCM_c405RdDBus[37]),
     .ISOCMC405RDDBUS38(           ISOCM_c405RdDBus[38]),
     .ISOCMC405RDDBUS39(           ISOCM_c405RdDBus[39]),
     .ISOCMC405RDDBUS40(           ISOCM_c405RdDBus[40]),
     .ISOCMC405RDDBUS41(           ISOCM_c405RdDBus[41]),
     .ISOCMC405RDDBUS42(           ISOCM_c405RdDBus[42]),
     .ISOCMC405RDDBUS43(           ISOCM_c405RdDBus[43]),
     .ISOCMC405RDDBUS44(           ISOCM_c405RdDBus[44]),
     .ISOCMC405RDDBUS45(           ISOCM_c405RdDBus[45]),
     .ISOCMC405RDDBUS46(           ISOCM_c405RdDBus[46]),
     .ISOCMC405RDDBUS47(           ISOCM_c405RdDBus[47]),
     .ISOCMC405RDDBUS48(           ISOCM_c405RdDBus[48]),
     .ISOCMC405RDDBUS49(           ISOCM_c405RdDBus[49]),
     .ISOCMC405RDDBUS50(           ISOCM_c405RdDBus[50]),
     .ISOCMC405RDDBUS51(           ISOCM_c405RdDBus[51]),
     .ISOCMC405RDDBUS52(           ISOCM_c405RdDBus[52]),
     .ISOCMC405RDDBUS53(           ISOCM_c405RdDBus[53]),
     .ISOCMC405RDDBUS54(           ISOCM_c405RdDBus[54]),
     .ISOCMC405RDDBUS55(           ISOCM_c405RdDBus[55]),
     .ISOCMC405RDDBUS56(           ISOCM_c405RdDBus[56]),
     .ISOCMC405RDDBUS57(           ISOCM_c405RdDBus[57]),
     .ISOCMC405RDDBUS58(           ISOCM_c405RdDBus[58]),
     .ISOCMC405RDDBUS59(           ISOCM_c405RdDBus[59]),
     .ISOCMC405RDDBUS60(           ISOCM_c405RdDBus[60]),
     .ISOCMC405RDDBUS61(           ISOCM_c405RdDBus[61]),
     .ISOCMC405RDDBUS62(           ISOCM_c405RdDBus[62]),
     .ISOCMC405RDDBUS63(           ISOCM_c405RdDBus[63]),
     .ISOCMC405RDDVALID0(          ISOCM_c405RdDValid[0]),
     .ISOCMC405RDDVALID1(          ISOCM_c405RdDValid[1]),
     .JTGC405BNDSCANTDO(           JTG_c405BndScanTDO),
     .JTGC405TCK(                  JTG_c405TCK),
     .JTGC405TDI(                  JTG_c405TDI),
     .JTGC405TMS(                  JTG_c405TMS),
     .JTGC405TRSTNEG(              JTG_c405TRST_NEG),
     .TESTC405BISTCCLK(            TEST_c405BistCClk),
     .TESTC405CNTLPOINT(           TEST_c405CntlPoint),
     .TESTC405TESTM1(              TEST_c405TestM1),
     .TESTC405TESTM3(              TEST_c405TestM3),
     .PLBC405DCUADDRACK(           PLB_c405DcuAddrAck),
     .PLBC405DCUBUSY(              PLB_c405DcuBusy),
     .PLBC405DCUERR(               PLB_c405DcuErr),
     .PLBC405DCURDDACK(            PLB_c405DcuRdDAck),
     .PLBC405DCURDDBUS00(          PLB_c405DcuRdDBus[0]),
     .PLBC405DCURDDBUS01(          PLB_c405DcuRdDBus[1]),
     .PLBC405DCURDDBUS02(          PLB_c405DcuRdDBus[2]),
     .PLBC405DCURDDBUS03(          PLB_c405DcuRdDBus[3]),
     .PLBC405DCURDDBUS04(          PLB_c405DcuRdDBus[4]),
     .PLBC405DCURDDBUS05(          PLB_c405DcuRdDBus[5]),
     .PLBC405DCURDDBUS06(          PLB_c405DcuRdDBus[6]),
     .PLBC405DCURDDBUS07(          PLB_c405DcuRdDBus[7]),
     .PLBC405DCURDDBUS08(          PLB_c405DcuRdDBus[8]),
     .PLBC405DCURDDBUS09(          PLB_c405DcuRdDBus[9]),
     .PLBC405DCURDDBUS10(          PLB_c405DcuRdDBus[10]),
     .PLBC405DCURDDBUS11(          PLB_c405DcuRdDBus[11]),
     .PLBC405DCURDDBUS12(          PLB_c405DcuRdDBus[12]),
     .PLBC405DCURDDBUS13(          PLB_c405DcuRdDBus[13]),
     .PLBC405DCURDDBUS14(          PLB_c405DcuRdDBus[14]),
     .PLBC405DCURDDBUS15(          PLB_c405DcuRdDBus[15]),
     .PLBC405DCURDDBUS16(          PLB_c405DcuRdDBus[16]),
     .PLBC405DCURDDBUS17(          PLB_c405DcuRdDBus[17]),
     .PLBC405DCURDDBUS18(          PLB_c405DcuRdDBus[18]),
     .PLBC405DCURDDBUS19(          PLB_c405DcuRdDBus[19]),
     .PLBC405DCURDDBUS20(          PLB_c405DcuRdDBus[20]),
     .PLBC405DCURDDBUS21(          PLB_c405DcuRdDBus[21]),
     .PLBC405DCURDDBUS22(          PLB_c405DcuRdDBus[22]),
     .PLBC405DCURDDBUS23(          PLB_c405DcuRdDBus[23]),
     .PLBC405DCURDDBUS24(          PLB_c405DcuRdDBus[24]),
     .PLBC405DCURDDBUS25(          PLB_c405DcuRdDBus[25]),
     .PLBC405DCURDDBUS26(          PLB_c405DcuRdDBus[26]),
     .PLBC405DCURDDBUS27(          PLB_c405DcuRdDBus[27]),
     .PLBC405DCURDDBUS28(          PLB_c405DcuRdDBus[28]),
     .PLBC405DCURDDBUS29(          PLB_c405DcuRdDBus[29]),
     .PLBC405DCURDDBUS30(          PLB_c405DcuRdDBus[30]),
     .PLBC405DCURDDBUS31(          PLB_c405DcuRdDBus[31]),
     .PLBC405DCURDDBUS32(          PLB_c405DcuRdDBus[32]),
     .PLBC405DCURDDBUS33(          PLB_c405DcuRdDBus[33]),
     .PLBC405DCURDDBUS34(          PLB_c405DcuRdDBus[34]),
     .PLBC405DCURDDBUS35(          PLB_c405DcuRdDBus[35]),
     .PLBC405DCURDDBUS36(          PLB_c405DcuRdDBus[36]),
     .PLBC405DCURDDBUS37(          PLB_c405DcuRdDBus[37]),
     .PLBC405DCURDDBUS38(          PLB_c405DcuRdDBus[38]),
     .PLBC405DCURDDBUS39(          PLB_c405DcuRdDBus[39]),
     .PLBC405DCURDDBUS40(          PLB_c405DcuRdDBus[40]),
     .PLBC405DCURDDBUS41(          PLB_c405DcuRdDBus[41]),
     .PLBC405DCURDDBUS42(          PLB_c405DcuRdDBus[42]),
     .PLBC405DCURDDBUS43(          PLB_c405DcuRdDBus[43]),
     .PLBC405DCURDDBUS44(          PLB_c405DcuRdDBus[44]),
     .PLBC405DCURDDBUS45(          PLB_c405DcuRdDBus[45]),
     .PLBC405DCURDDBUS46(          PLB_c405DcuRdDBus[46]),
     .PLBC405DCURDDBUS47(          PLB_c405DcuRdDBus[47]),
     .PLBC405DCURDDBUS48(          PLB_c405DcuRdDBus[48]),
     .PLBC405DCURDDBUS49(          PLB_c405DcuRdDBus[49]),
     .PLBC405DCURDDBUS50(          PLB_c405DcuRdDBus[50]),
     .PLBC405DCURDDBUS51(          PLB_c405DcuRdDBus[51]),
     .PLBC405DCURDDBUS52(          PLB_c405DcuRdDBus[52]),
     .PLBC405DCURDDBUS53(          PLB_c405DcuRdDBus[53]),
     .PLBC405DCURDDBUS54(          PLB_c405DcuRdDBus[54]),
     .PLBC405DCURDDBUS55(          PLB_c405DcuRdDBus[55]),
     .PLBC405DCURDDBUS56(          PLB_c405DcuRdDBus[56]),
     .PLBC405DCURDDBUS57(          PLB_c405DcuRdDBus[57]),
     .PLBC405DCURDDBUS58(          PLB_c405DcuRdDBus[58]),
     .PLBC405DCURDDBUS59(          PLB_c405DcuRdDBus[59]),
     .PLBC405DCURDDBUS60(          PLB_c405DcuRdDBus[60]),
     .PLBC405DCURDDBUS61(          PLB_c405DcuRdDBus[61]),
     .PLBC405DCURDDBUS62(          PLB_c405DcuRdDBus[62]),
     .PLBC405DCURDDBUS63(          PLB_c405DcuRdDBus[63]),
     .PLBC405DCURDWDADDR1(         PLB_c405DcuRdWdAddr[1]),
     .PLBC405DCURDWDADDR2(         PLB_c405DcuRdWdAddr[2]),
     .PLBC405DCURDWDADDR3(         PLB_c405DcuRdWdAddr[3]),
     .PLBC405DCUSSIZE1(            PLB_c405DcuSSize1),
     .PLBC405DCUWRDACK(            PLB_c405DcuWrDAck),
     .PLBC405ICUADDRACK(           PLB_c405IcuAddrAck),
     .PLBC405ICUBUSY(              PLB_c405IcuBusy),
     .PLBC405ICUERR(               PLB_c405IcuErr),
     .PLBC405ICURDDACK(            PLB_c405IcuRdDAck),
     .PLBC405ICURDDBUS00(          PLB_c405IcuRdDBus[0]),
     .PLBC405ICURDDBUS01(          PLB_c405IcuRdDBus[1]),
     .PLBC405ICURDDBUS02(          PLB_c405IcuRdDBus[2]),
     .PLBC405ICURDDBUS03(          PLB_c405IcuRdDBus[3]),
     .PLBC405ICURDDBUS04(          PLB_c405IcuRdDBus[4]),
     .PLBC405ICURDDBUS05(          PLB_c405IcuRdDBus[5]),
     .PLBC405ICURDDBUS06(          PLB_c405IcuRdDBus[6]),
     .PLBC405ICURDDBUS07(          PLB_c405IcuRdDBus[7]),
     .PLBC405ICURDDBUS08(          PLB_c405IcuRdDBus[8]),
     .PLBC405ICURDDBUS09(          PLB_c405IcuRdDBus[9]),
     .PLBC405ICURDDBUS10(          PLB_c405IcuRdDBus[10]),
     .PLBC405ICURDDBUS11(          PLB_c405IcuRdDBus[11]),
     .PLBC405ICURDDBUS12(          PLB_c405IcuRdDBus[12]),
     .PLBC405ICURDDBUS13(          PLB_c405IcuRdDBus[13]),
     .PLBC405ICURDDBUS14(          PLB_c405IcuRdDBus[14]),
     .PLBC405ICURDDBUS15(          PLB_c405IcuRdDBus[15]),
     .PLBC405ICURDDBUS16(          PLB_c405IcuRdDBus[16]),
     .PLBC405ICURDDBUS17(          PLB_c405IcuRdDBus[17]),
     .PLBC405ICURDDBUS18(          PLB_c405IcuRdDBus[18]),
     .PLBC405ICURDDBUS19(          PLB_c405IcuRdDBus[19]),
     .PLBC405ICURDDBUS20(          PLB_c405IcuRdDBus[20]),
     .PLBC405ICURDDBUS21(          PLB_c405IcuRdDBus[21]),
     .PLBC405ICURDDBUS22(          PLB_c405IcuRdDBus[22]),
     .PLBC405ICURDDBUS23(          PLB_c405IcuRdDBus[23]),
     .PLBC405ICURDDBUS24(          PLB_c405IcuRdDBus[24]),
     .PLBC405ICURDDBUS25(          PLB_c405IcuRdDBus[25]),
     .PLBC405ICURDDBUS26(          PLB_c405IcuRdDBus[26]),
     .PLBC405ICURDDBUS27(          PLB_c405IcuRdDBus[27]),
     .PLBC405ICURDDBUS28(          PLB_c405IcuRdDBus[28]),
     .PLBC405ICURDDBUS29(          PLB_c405IcuRdDBus[29]),
     .PLBC405ICURDDBUS30(          PLB_c405IcuRdDBus[30]),
     .PLBC405ICURDDBUS31(          PLB_c405IcuRdDBus[31]),
     .PLBC405ICURDDBUS32(          PLB_c405IcuRdDBus[32]),
     .PLBC405ICURDDBUS33(          PLB_c405IcuRdDBus[33]),
     .PLBC405ICURDDBUS34(          PLB_c405IcuRdDBus[34]),
     .PLBC405ICURDDBUS35(          PLB_c405IcuRdDBus[35]),
     .PLBC405ICURDDBUS36(          PLB_c405IcuRdDBus[36]),
     .PLBC405ICURDDBUS37(          PLB_c405IcuRdDBus[37]),
     .PLBC405ICURDDBUS38(          PLB_c405IcuRdDBus[38]),
     .PLBC405ICURDDBUS39(          PLB_c405IcuRdDBus[39]),
     .PLBC405ICURDDBUS40(          PLB_c405IcuRdDBus[40]),
     .PLBC405ICURDDBUS41(          PLB_c405IcuRdDBus[41]),
     .PLBC405ICURDDBUS42(          PLB_c405IcuRdDBus[42]),
     .PLBC405ICURDDBUS43(          PLB_c405IcuRdDBus[43]),
     .PLBC405ICURDDBUS44(          PLB_c405IcuRdDBus[44]),
     .PLBC405ICURDDBUS45(          PLB_c405IcuRdDBus[45]),
     .PLBC405ICURDDBUS46(          PLB_c405IcuRdDBus[46]),
     .PLBC405ICURDDBUS47(          PLB_c405IcuRdDBus[47]),
     .PLBC405ICURDDBUS48(          PLB_c405IcuRdDBus[48]),
     .PLBC405ICURDDBUS49(          PLB_c405IcuRdDBus[49]),
     .PLBC405ICURDDBUS50(          PLB_c405IcuRdDBus[50]),
     .PLBC405ICURDDBUS51(          PLB_c405IcuRdDBus[51]),
     .PLBC405ICURDDBUS52(          PLB_c405IcuRdDBus[52]),
     .PLBC405ICURDDBUS53(          PLB_c405IcuRdDBus[53]),
     .PLBC405ICURDDBUS54(          PLB_c405IcuRdDBus[54]),
     .PLBC405ICURDDBUS55(          PLB_c405IcuRdDBus[55]),
     .PLBC405ICURDDBUS56(          PLB_c405IcuRdDBus[56]),
     .PLBC405ICURDDBUS57(          PLB_c405IcuRdDBus[57]),
     .PLBC405ICURDDBUS58(          PLB_c405IcuRdDBus[58]),
     .PLBC405ICURDDBUS59(          PLB_c405IcuRdDBus[59]),
     .PLBC405ICURDDBUS60(          PLB_c405IcuRdDBus[60]),
     .PLBC405ICURDDBUS61(          PLB_c405IcuRdDBus[61]),
     .PLBC405ICURDDBUS62(          PLB_c405IcuRdDBus[62]),
     .PLBC405ICURDDBUS63(          PLB_c405IcuRdDBus[63]),
     .PLBC405ICURDWDADDR1(         PLB_c405IcuRdWdAddr[1]),
     .PLBC405ICURDWDADDR2(         PLB_c405IcuRdWdAddr[2]),
     .PLBC405ICURDWDADDR3(         PLB_c405IcuRdWdAddr[3]),
     .PLBC405ICUSSIZE1(            PLB_c405IcuSSize1),
     .RSTC405RESETCHIP(            RST_c405ResetChip),
     .RSTC405RESETCORE(            RST_c405ResetCore),
     .RSTC405RESETSYSTEM(          RST_c405ResetSystem),
     .TIEC405APUDIVEN(             TIE_c405ApuDivEn),
     .TIEC405APUPRESENT(           TIE_c405ApuPresent),
     .TIEC405DETERMINISTICMULT(    TIE_c405DeterministicMult),
     .TIEC405DISOPERANDFWD(        TIE_c405DisOperandFwd),
     .TIEC405MMUEN(                TIE_c405MmuEn),
     .TIEC405PVR00(                TIE_c405PVR[0]),
     .TIEC405PVR01(                TIE_c405PVR[1]),
     .TIEC405PVR02(                TIE_c405PVR[2]),
     .TIEC405PVR03(                TIE_c405PVR[3]),
     .TIEC405PVR04(                TIE_c405PVR[4]),
     .TIEC405PVR05(                TIE_c405PVR[5]),
     .TIEC405PVR06(                TIE_c405PVR[6]),
     .TIEC405PVR07(                TIE_c405PVR[7]),
     .TIEC405PVR08(                TIE_c405PVR[8]),
     .TIEC405PVR09(                TIE_c405PVR[9]),
     .TIEC405PVR10(                TIE_c405PVR[10]),
     .TIEC405PVR11(                TIE_c405PVR[11]),
     .TIEC405PVR12(                TIE_c405PVR[12]),
     .TIEC405PVR13(                TIE_c405PVR[13]),
     .TIEC405PVR14(                TIE_c405PVR[14]),
     .TIEC405PVR15(                TIE_c405PVR[15]),
     .TIEC405PVR16(                TIE_c405PVR[16]),
     .TIEC405PVR17(                TIE_c405PVR[17]),
     .TIEC405PVR18(                TIE_c405PVR[18]),
     .TIEC405PVR19(                TIE_c405PVR[19]),
     .TIEC405PVR20(                TIE_c405PVR[20]),
     .TIEC405PVR21(                TIE_c405PVR[21]),
     .TIEC405PVR22(                TIE_c405PVR[22]),
     .TIEC405PVR23(                TIE_c405PVR[23]),
     .TIEC405PVR24(                TIE_c405PVR[24]),
     .TIEC405PVR25(                TIE_c405PVR[25]),
     .TIEC405PVR26(                TIE_c405PVR[26]),
     .TIEC405PVR27(                TIE_c405PVR[27]),
     .TIEC405PVR28(                TIE_c405PVR[28]),
     .TIEC405PVR29(                TIE_c405PVR[29]),
     .TIEC405PVR30(                TIE_c405PVR[30]),
     .TIEC405PVR31(                TIE_c405PVR[31]),
     .TRCC405TRACEDISABLE(         TRC_c405TraceDisable),
     .TRCC405TRIGGEREVENTIN(       TRC_c405TriggerEventIn),
     .C405BISTPEPSPF00(            C405_bistPepsPF[0]),
     .C405BISTPEPSPF01(            C405_bistPepsPF[1]),
     .C405BISTPEPSPF02(            C405_bistPepsPF[2]),
     .TESTC405CE0EVS(              TEST_c405CE0EVS),
     .TESTC405BISTCE0STCLK(        TEST_c405BistCE0StClk),
     .TESTC405BISTCE1ENABLE(       TEST_c405BistCE1Enable),
     .TESTC405BISTCE1MODE(         TEST_c405BistCE1Mode),
     .CPMC405PLBSYNCCLOCK(         CPM_c405PlbSyncClock),
     .CPMC405SYNCBYPASS(           CPM_c405SyncBypass),
     .TIEC405CLOCKENABLE(          TIE_c405ClockEnable),
     .TIEC405DUTYENABLE(           TIE_c405DutyEnable),
     .CPMC405PLBSAMPLECYCLEALT(    CPM_c405PlbSampleCycleAlt),

     .C405TESTSCANOUT0   ( C405_testScanOut[0]),
     .C405TESTSCANOUT1   ( C405_testScanOut[1]),
     .C405TESTSCANOUT2   ( C405_testScanOut[2]),
     .C405TESTSCANOUT3   ( C405_testScanOut[3]),
     .C405TESTSCANOUT4   ( C405_testScanOut[4]),
     .C405TESTSCANOUT5   ( C405_testScanOut[5]),
     .C405TESTSCANOUT6   ( C405_testScanOut[6]),
     .C405TESTSCANOUT7   ( C405_testScanOut[7]),
     
     .TESTC405SCANIN0   ( TEST_c405ScanIn[0]),
     .TESTC405SCANIN1   ( TEST_c405ScanIn[1]),
     .TESTC405SCANIN2   ( TEST_c405ScanIn[2]),
     .TESTC405SCANIN3   ( TEST_c405ScanIn[3]),
     .TESTC405SCANIN4   ( TEST_c405ScanIn[4]),
     .TESTC405SCANIN5   ( TEST_c405ScanIn[5]),
     .TESTC405SCANIN6   ( TEST_c405ScanIn[6]),
     .TESTC405SCANIN7   ( TEST_c405ScanIn[7]),
     .TESTC405SCANENABLE (TEST_c405ScanEnable),
     .TESTC405TESTMODE (TEST_c405TestMode),

     .BISTC405DCUBISTDEBUGSI00   ( BIST_c405dcuBistDebugSi[0]),
     .BISTC405DCUBISTDEBUGSI01   ( BIST_c405dcuBistDebugSi[1]),
     .BISTC405DCUBISTDEBUGSI02   ( BIST_c405dcuBistDebugSi[2]),
     .BISTC405DCUBISTDEBUGSI03   ( BIST_c405dcuBistDebugSi[3]),
     .C405BISTDCUBISTDEBUGSO00   ( C405_bistdcuBistDebugSo[0]),
     .C405BISTDCUBISTDEBUGSO01   ( C405_bistdcuBistDebugSo[1]),
     .C405BISTDCUBISTDEBUGSO02   ( C405_bistdcuBistDebugSo[2]),
     .C405BISTDCUBISTDEBUGSO03   ( C405_bistdcuBistDebugSo[3]),
     .BISTC405DCUBISTDEBUGEN00   ( BIST_c405dcuBistDebugEn[0]),
     .BISTC405DCUBISTDEBUGEN01   ( BIST_c405dcuBistDebugEn[1]),
     .BISTC405DCUBISTDEBUGEN02   ( BIST_c405dcuBistDebugEn[2]),
     .BISTC405DCUBISTDEBUGEN03   ( BIST_c405dcuBistDebugEn[3]),
     .BISTC405DCUBISTMODEREGIN00   ( BIST_c405dcuBistModeRegIn[0]),
     .BISTC405DCUBISTMODEREGIN01   ( BIST_c405dcuBistModeRegIn[1]),
     .BISTC405DCUBISTMODEREGIN02   ( BIST_c405dcuBistModeRegIn[2]),
     .BISTC405DCUBISTMODEREGIN03   ( BIST_c405dcuBistModeRegIn[3]),
     .BISTC405DCUBISTMODEREGIN04   ( BIST_c405dcuBistModeRegIn[4]),
     .BISTC405DCUBISTMODEREGIN05   ( BIST_c405dcuBistModeRegIn[5]),
     .BISTC405DCUBISTMODEREGIN06   ( BIST_c405dcuBistModeRegIn[6]),
     .BISTC405DCUBISTMODEREGIN07   ( BIST_c405dcuBistModeRegIn[7]),
     .BISTC405DCUBISTMODEREGIN08   ( BIST_c405dcuBistModeRegIn[8]),
     .BISTC405DCUBISTMODEREGIN09   ( BIST_c405dcuBistModeRegIn[9]),
     .BISTC405DCUBISTMODEREGIN10   ( BIST_c405dcuBistModeRegIn[10]),
     .BISTC405DCUBISTMODEREGIN11   ( BIST_c405dcuBistModeRegIn[11]),
     .BISTC405DCUBISTMODEREGIN12   ( BIST_c405dcuBistModeRegIn[12]),
     .BISTC405DCUBISTMODEREGIN13   ( BIST_c405dcuBistModeRegIn[13]),
     .BISTC405DCUBISTMODEREGIN14   ( BIST_c405dcuBistModeRegIn[14]),
     .BISTC405DCUBISTMODEREGIN15   ( BIST_c405dcuBistModeRegIn[15]),
     .BISTC405DCUBISTMODEREGIN16   ( BIST_c405dcuBistModeRegIn[16]),
     .BISTC405DCUBISTMODEREGIN17   ( BIST_c405dcuBistModeRegIn[17]),
     .BISTC405DCUBISTMODEREGIN18   ( BIST_c405dcuBistModeRegIn[18]),
     .C405BISTDCUBISTMODEREGOUT00   ( C405_bistdcuBistModeRegOut[0]),
     .C405BISTDCUBISTMODEREGOUT01   ( C405_bistdcuBistModeRegOut[1]),
     .C405BISTDCUBISTMODEREGOUT02   ( C405_bistdcuBistModeRegOut[2]),
     .C405BISTDCUBISTMODEREGOUT03   ( C405_bistdcuBistModeRegOut[3]),
     .C405BISTDCUBISTMODEREGOUT04   ( C405_bistdcuBistModeRegOut[4]),
     .C405BISTDCUBISTMODEREGOUT05   ( C405_bistdcuBistModeRegOut[5]),
     .C405BISTDCUBISTMODEREGOUT06   ( C405_bistdcuBistModeRegOut[6]),
     .C405BISTDCUBISTMODEREGOUT07   ( C405_bistdcuBistModeRegOut[7]),
     .C405BISTDCUBISTMODEREGOUT08   ( C405_bistdcuBistModeRegOut[8]),
     .C405BISTDCUBISTMODEREGOUT09   ( C405_bistdcuBistModeRegOut[9]),
     .C405BISTDCUBISTMODEREGOUT10   ( C405_bistdcuBistModeRegOut[10]),
     .C405BISTDCUBISTMODEREGOUT11   ( C405_bistdcuBistModeRegOut[11]),
     .C405BISTDCUBISTMODEREGOUT12   ( C405_bistdcuBistModeRegOut[12]),
     .C405BISTDCUBISTMODEREGOUT13   ( C405_bistdcuBistModeRegOut[13]),
     .C405BISTDCUBISTMODEREGOUT14   ( C405_bistdcuBistModeRegOut[14]),
     .C405BISTDCUBISTMODEREGOUT15   ( C405_bistdcuBistModeRegOut[15]),
     .C405BISTDCUBISTMODEREGOUT16   ( C405_bistdcuBistModeRegOut[16]),
     .C405BISTDCUBISTMODEREGOUT17   ( C405_bistdcuBistModeRegOut[17]),
     .C405BISTDCUBISTMODEREGOUT18   ( C405_bistdcuBistModeRegOut[18]),
     .BISTC405DCUBISTPARALLELDR   ( BIST_c405dcuBistParallelDr),
     .BISTC405DCUBISTMODEREGSI   ( BIST_c405dcuBistModeRegSi),
     .C405BISTDCUBISTMODEREGSO   ( C405_bistdcuBistModeRegSo),
     .BISTC405DCUBISTSHIFTDR   ( BIST_c405dcuBistShiftDr),
     .BISTC405DCUBISTMBRUN   ( BIST_c405dcuBistMbRun),

     .BISTC405ICUBISTDEBUGSI00   ( BIST_c405icuBistDebugSi[0]),
     .BISTC405ICUBISTDEBUGSI01   ( BIST_c405icuBistDebugSi[1]),
     .BISTC405ICUBISTDEBUGSI02   ( BIST_c405icuBistDebugSi[2]),
     .BISTC405ICUBISTDEBUGSI03   ( BIST_c405icuBistDebugSi[3]),
     .C405BISTICUBISTDEBUGSO00   ( C405_bisticuBistDebugSo[0]),
     .C405BISTICUBISTDEBUGSO01   ( C405_bisticuBistDebugSo[1]),
     .C405BISTICUBISTDEBUGSO02   ( C405_bisticuBistDebugSo[2]),
     .C405BISTICUBISTDEBUGSO03   ( C405_bisticuBistDebugSo[3]),
     .BISTC405ICUBISTDEBUGEN00   ( BIST_c405icuBistDebugEn[0]),
     .BISTC405ICUBISTDEBUGEN01   ( BIST_c405icuBistDebugEn[1]),
     .BISTC405ICUBISTDEBUGEN02   ( BIST_c405icuBistDebugEn[2]),
     .BISTC405ICUBISTDEBUGEN03   ( BIST_c405icuBistDebugEn[3]),
     .BISTC405ICUBISTMODEREGIN00   ( BIST_c405icuBistModeRegIn[0]),
     .BISTC405ICUBISTMODEREGIN01   ( BIST_c405icuBistModeRegIn[1]),
     .BISTC405ICUBISTMODEREGIN02   ( BIST_c405icuBistModeRegIn[2]),
     .BISTC405ICUBISTMODEREGIN03   ( BIST_c405icuBistModeRegIn[3]),
     .BISTC405ICUBISTMODEREGIN04   ( BIST_c405icuBistModeRegIn[4]),
     .BISTC405ICUBISTMODEREGIN05   ( BIST_c405icuBistModeRegIn[5]),
     .BISTC405ICUBISTMODEREGIN06   ( BIST_c405icuBistModeRegIn[6]),
     .BISTC405ICUBISTMODEREGIN07   ( BIST_c405icuBistModeRegIn[7]),
     .BISTC405ICUBISTMODEREGIN08   ( BIST_c405icuBistModeRegIn[8]),
     .BISTC405ICUBISTMODEREGIN09   ( BIST_c405icuBistModeRegIn[9]),
     .BISTC405ICUBISTMODEREGIN10   ( BIST_c405icuBistModeRegIn[10]),
     .BISTC405ICUBISTMODEREGIN11   ( BIST_c405icuBistModeRegIn[11]),
     .BISTC405ICUBISTMODEREGIN12   ( BIST_c405icuBistModeRegIn[12]),
     .BISTC405ICUBISTMODEREGIN13   ( BIST_c405icuBistModeRegIn[13]),
     .BISTC405ICUBISTMODEREGIN14   ( BIST_c405icuBistModeRegIn[14]),
     .BISTC405ICUBISTMODEREGIN15   ( BIST_c405icuBistModeRegIn[15]),
     .BISTC405ICUBISTMODEREGIN16   ( BIST_c405icuBistModeRegIn[16]),
     .BISTC405ICUBISTMODEREGIN17   ( BIST_c405icuBistModeRegIn[17]),
     .BISTC405ICUBISTMODEREGIN18   ( BIST_c405icuBistModeRegIn[18]),
     .C405BISTICUBISTMODEREGOUT00   ( C405_bisticuBistModeRegOut[0]),
     .C405BISTICUBISTMODEREGOUT01   ( C405_bisticuBistModeRegOut[1]),
     .C405BISTICUBISTMODEREGOUT02   ( C405_bisticuBistModeRegOut[2]),
     .C405BISTICUBISTMODEREGOUT03   ( C405_bisticuBistModeRegOut[3]),
     .C405BISTICUBISTMODEREGOUT04   ( C405_bisticuBistModeRegOut[4]),
     .C405BISTICUBISTMODEREGOUT05   ( C405_bisticuBistModeRegOut[5]),
     .C405BISTICUBISTMODEREGOUT06   ( C405_bisticuBistModeRegOut[6]),
     .C405BISTICUBISTMODEREGOUT07   ( C405_bisticuBistModeRegOut[7]),
     .C405BISTICUBISTMODEREGOUT08   ( C405_bisticuBistModeRegOut[8]),
     .C405BISTICUBISTMODEREGOUT09   ( C405_bisticuBistModeRegOut[9]),
     .C405BISTICUBISTMODEREGOUT10   ( C405_bisticuBistModeRegOut[10]),
     .C405BISTICUBISTMODEREGOUT11   ( C405_bisticuBistModeRegOut[11]),
     .C405BISTICUBISTMODEREGOUT12   ( C405_bisticuBistModeRegOut[12]),
     .C405BISTICUBISTMODEREGOUT13   ( C405_bisticuBistModeRegOut[13]),
     .C405BISTICUBISTMODEREGOUT14   ( C405_bisticuBistModeRegOut[14]),
     .C405BISTICUBISTMODEREGOUT15   ( C405_bisticuBistModeRegOut[15]),
     .C405BISTICUBISTMODEREGOUT16   ( C405_bisticuBistModeRegOut[16]),
     .C405BISTICUBISTMODEREGOUT17   ( C405_bisticuBistModeRegOut[17]),
     .C405BISTICUBISTMODEREGOUT18   ( C405_bisticuBistModeRegOut[18]),
     .BISTC405ICUBISTPARALLELDR   ( BIST_c405icuBistParallelDr),
     .BISTC405ICUBISTMODEREGSI   ( BIST_c405icuBistModeRegSi),
     .C405BISTICUBISTMODEREGSO   ( C405_bisticuBistModeRegSo),
     .BISTC405ICUBISTSHIFTDR   ( BIST_c405icuBistShiftDr),
     .BISTC405ICUBISTMBRUN   ( BIST_c405icuBistMbRun)
//      .BISTC405ICUBISTDEBUGSI   ( BIST_c405icuBistDebugSi),
//      .C405BISTICUBISTDEBUGSO   ( C405_bisticuBistDebugSo),
//      .BISTC405ICUBISTDEBUGEN   ( BIST_c405icuBistDebugEn),
//      .BISTC405ICUBISTMODEREGIN   ( BIST_c405icuBistModeRegIn),
//      .C405BISTICUBISTMODEREGOUT   ( C405_bisticuBistModeRegOut),
//      .BISTC405ICUBISTPARALLELDR   ( BIST_c405icuBistParallelDr),
//      .BISTC405ICUBISTMODEREGSI   ( BIST_c405icuBistModeRegSi),
//      .C405BISTICUBISTMODEREGSO   ( C405_bisticuBistModeRegSo),
//      .BISTC405ICUBISTSHIFTDR   ( BIST_c405icuBistShiftDr),
//      .BISTC405ICUBISTMBRUN   ( BIST_c405icuBistMbRun)

     );

endmodule
