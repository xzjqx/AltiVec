library verilog;
use verilog.vl_types.all;
entity p405s_test_top is
    generic(
        simulation_cycle: integer := 10
    );
end p405s_test_top;
