library verilog;
use verilog.vl_types.all;
entity p405s_pipeCntl is
    port(
        PCL_dcdAregLoadUse: out    vl_logic;
        PCL_aPortRregBypass: out    vl_logic;
        PCL_abRegE1     : out    vl_logic;
        PCL_aRegE2      : out    vl_logic;
        PCL_dcdBregLoadUse: out    vl_logic;
        PCL_bPortRregBypass: out    vl_logic;
        PCL_bRegE2      : out    vl_logic;
        PCL_blkFlush    : out    vl_logic;
        PCL_dRegBypassMuxSel: out    vl_logic;
        PCL_dRegE1      : out    vl_logic;
        PCL_dcdHoldForIfb: out    vl_logic_vector(0 to 2);
        PCL_dofDRegE1   : out    vl_logic;
        PCL_dofDRegMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exeIarHold  : out    vl_logic;
        PCL_mfDCR       : out    vl_logic;
        PCL_mtDCR       : out    vl_logic;
        PCL_gateZeroToAreg: out    vl_logic;
        PCL_gateZeroToSreg: out    vl_logic;
        PCL_holdCIn     : out    vl_logic;
        PCL_ldAdjE1     : out    vl_logic;
        PCL_ldAdjMuxSel : out    vl_logic_vector(0 to 1);
        PCL_ldMuxSel    : out    vl_logic_vector(0 to 7);
        PCL_lwbLpWrEn   : out    vl_logic;
        PCL_resultRegE1 : out    vl_logic;
        PCL_resultRegE2 : out    vl_logic;
        PCL_dcdSregLoadUse: out    vl_logic;
        PCL_sPortRregBypass: out    vl_logic;
        PCL_sRegE1      : out    vl_logic;
        PCL_sRegE2      : out    vl_logic;
        PCL_sraRegE1    : out    vl_logic;
        PCL_dIcmpForStep: out    vl_logic;
        PCL_srmRegE1    : out    vl_logic;
        PCL_srmRegE2    : out    vl_logic_vector(0 to 2);
        PCL_wbHold      : out    vl_logic;
        PCL_xerL2Hold   : out    vl_logic;
        countE2         : out    vl_logic;
        dcdStringImmediate: out    vl_logic;
        dcdXerTBCUpdInstr: out    vl_logic;
        exeClearOrFlush : out    vl_logic;
        exeE1           : out    vl_logic;
        exeE2           : out    vl_logic;
        exeLpAddrE2     : out    vl_logic;
        exeLpMuxSel     : out    vl_logic;
        exeRpAddrE2     : out    vl_logic;
        gtErr           : out    vl_logic;
        loadSteerMuxSel : out    vl_logic;
        lwbE1           : out    vl_logic;
        nxtWbLpWrEn     : out    vl_logic;
        storageStMachE2 : out    vl_logic;
        storeRSE2       : out    vl_logic;
        PCL_wbClearOrFlush: out    vl_logic;
        wbE1            : out    vl_logic;
        wbE2            : out    vl_logic;
        APU_exeBlkingMco: in     vl_logic;
        APU_exeBusy     : in     vl_logic;
        APU_exeNonBlkingMco: in     vl_logic;
        CB              : in     vl_logic;
        DCU_CA          : in     vl_logic;
        DCU_DA          : in     vl_logic;
        DCU_DOF         : in     vl_logic;
        EXE_admMco      : in     vl_logic;
        ICU_dsCA        : in     vl_logic;
        IFB_dcdFull     : in     vl_logic;
        gprLpeqRp       : in     vl_logic;
        MMU_BMCO        : in     vl_logic;
        MMU_wbHold      : in     vl_logic;
        NplaApRdEn      : in     vl_logic;
        NplaAregEn      : in     vl_logic;
        NplaBpRdEn      : in     vl_logic;
        NplaBregEn      : in     vl_logic;
        plaSpRdEn       : in     vl_logic;
        NplaSregEn      : in     vl_logic;
        OCM_dsComplete  : in     vl_logic;
        OCM_DOF         : in     vl_logic;
        VCT_exeSuppress : in     vl_logic;
        VCT_wbFlush     : in     vl_logic;
        coreReset       : in     vl_logic;
        dcdRAL2         : in     vl_logic_vector(0 to 4);
        dcdSPRN         : in     vl_logic_vector(0 to 9);
        XXX_dcrAck      : in     vl_logic;
        exeEaCalc       : in     vl_logic;
        exeLSSMIURA     : in     vl_logic_vector(0 to 5);
        lwbLpEqdcdApAddr: in     vl_logic;
        lwbLpEqdcdBpAddr: in     vl_logic;
        lwbLpEqdcdSpAddr: in     vl_logic;
        exeMfdcr        : in     vl_logic;
        exeMtdcr        : in     vl_logic;
        exeRTeqRA       : in     vl_logic;
        exeRTeqRB       : in     vl_logic;
        exeRpEqdcdApAddr: in     vl_logic;
        exeRpEqdcdBpAddr: in     vl_logic;
        exeRpEqdcdSpAddr: in     vl_logic;
        exeRpEqlwbLpAddr: in     vl_logic;
        exeRpEqwbLpAddr : in     vl_logic;
        exeRpWrEn       : in     vl_logic;
        exeStrgSt       : in     vl_logic_vector(0 to 2);
        ldAdjSel        : in     vl_logic_vector(1 to 3);
        lwbLpEqexeApAddr: in     vl_logic;
        lwbLpEqexeBpAddr: in     vl_logic;
        lwbLpEqexeSpAddr: in     vl_logic;
        nopStringIndexed: in     vl_logic;
        plaLSSMIURA     : in     vl_logic_vector(0 to 4);
        plaLogicalCntl  : in     vl_logic_vector(6 to 7);
        plaMtspr        : in     vl_logic;
        plaRaEq0Ck      : in     vl_logic;
        plaSrmEn        : in     vl_logic;
        priOp           : in     vl_logic_vector(0 to 5);
        strgEnd         : in     vl_logic;
        strgLpWrEn      : in     vl_logic;
        wbFull          : in     vl_logic;
        wbLoad          : in     vl_logic;
        wbLpEqdcdApAddr : in     vl_logic;
        wbLpEqdcdBpAddr : in     vl_logic;
        wbLpEqdcdSpAddr : in     vl_logic;
        wbLpWrEn        : in     vl_logic;
        sPortSelInc     : in     vl_logic;
        sprHold         : out    vl_logic;
        exeRpWrEnQ      : out    vl_logic;
        nxtExeFull      : out    vl_logic;
        exeFull         : in     vl_logic;
        IFB_exeCorrect  : in     vl_logic;
        IFB_trcPipeHold : in     vl_logic;
        wbRpAddrE2      : out    vl_logic;
        plaLpWrEn       : in     vl_logic;
        PCL_wbRpWrEn    : in     vl_logic;
        wbStrgLS        : in     vl_logic;
        PCL_exeAbort    : out    vl_logic;
        exeStwcx        : in     vl_logic;
        wbLwarx         : in     vl_logic;
        wbStwcx         : in     vl_logic;
        VCT_wbSuppress  : in     vl_logic;
        wbLpEqexeApAddr : in     vl_logic;
        wbLpEqexeBpAddr : in     vl_logic;
        wbLpEqexeSpAddr : in     vl_logic;
        exeApRdEn       : in     vl_logic;
        exeBpRdEn       : in     vl_logic;
        exeSpRdEn       : in     vl_logic;
        exeSpAddrE2     : out    vl_logic;
        PCL_exeAregLoadUse: out    vl_logic;
        PCL_exeBregLoadUse: out    vl_logic;
        PCL_exeSregLoadUse: out    vl_logic;
        EXE_divMco      : in     vl_logic;
        IFB_dcdBubble   : in     vl_logic;
        plaTrap         : in     vl_logic;
        exeSrmUnitEn    : in     vl_logic;
        NdcdApRdEn      : out    vl_logic;
        DCU_pclOcmLdPendNoWait: in     vl_logic;
        PCL_Rbit        : out    vl_logic;
        ICU_LDBE        : in     vl_logic;
        PCL_apuLwbLoadDV: out    vl_logic;
        PCL_apuTrcLoadEn: out    vl_logic;
        wbApuFpuLoad    : in     vl_logic;
        exeApuFpuOp     : in     vl_logic;
        IFB_exeFlush    : in     vl_logic;
        plaDcuOp        : in     vl_logic_vector(4 to 5);
        VCT_errorSprSuppress: in     vl_logic;
        DCU_firstCycCarStXltV: in     vl_logic;
        DBG_dvcRdEn     : in     vl_logic;
        DBG_dvcWrEn     : in     vl_logic;
        exeDcbz         : in     vl_logic;
        exeDcba         : in     vl_logic;
        exeMultEn       : in     vl_logic;
        exeDivEn        : in     vl_logic;
        exeMacEn        : in     vl_logic;
        PCL_apuExeHold  : out    vl_logic;
        PCL_apuExeFlush : out    vl_logic;
        EXE_trap        : in     vl_logic;
        PCL_exeTrap     : out    vl_logic;
        exe2Full        : in     vl_logic;
        plaMacEn        : in     vl_logic;
        DBG_icmpEn      : in     vl_logic;
        PCL_exeDvcHold  : out    vl_logic;
        PCL_wbStorageOp : in     vl_logic;
        PCL_exe2Hold    : out    vl_logic;
        EXE_multMco     : in     vl_logic;
        PCL_dvcCmpEn    : out    vl_logic;
        PCL_exe2IarE1   : out    vl_logic;
        PCL_exe2IarE2   : out    vl_logic;
        PCL_exe2DataE1  : out    vl_logic;
        PCL_exe2DataE2  : out    vl_logic;
        PCL_exe2ClearOrFlush: out    vl_logic;
        wbLdOrStWUD     : in     vl_logic;
        exeMacOrMultRpAddrE2: out    vl_logic;
        exeRpAddrMuxSel : out    vl_logic;
        dcdMmuSprDcd    : out    vl_logic_vector(0 to 8);
        PCL_trcLoadDV   : out    vl_logic;
        wbStrgC1        : in     vl_logic;
        PCL_wbDbgIcmp   : out    vl_logic;
        MMU_dsStatus    : in     vl_logic_vector(0 to 4);
        IFB_exeRfciL2   : in     vl_logic;
        IFB_exeRfiL2    : in     vl_logic;
        IFB_exeScL2     : in     vl_logic;
        VCT_wbFlushAsync: in     vl_logic;
        IFB_stepStL2    : in     vl_logic;
        PCL_mfDCRL2     : out    vl_logic;
        PCL_wbHoldNonErr: out    vl_logic;
        PCL_wbFullForPO : out    vl_logic;
        PCL_wbComplete  : out    vl_logic;
        PCL_apuDcdHold  : out    vl_logic;
        exeMorMRpEqdcdApAddr: in     vl_logic;
        exeMorMRpEqdcdBpAddr: in     vl_logic;
        lwbFullL2       : out    vl_logic;
        VCT_wbLoadSuppress: in     vl_logic;
        plaMultEn       : in     vl_logic;
        plaLogicalUnitEn: in     vl_logic;
        plaVal          : in     vl_logic;
        blkExeSpAddr    : in     vl_logic;
        storageStMachE1 : out    vl_logic;
        wbLpAddrE1      : out    vl_logic;
        PCL_exeHoldForCr: out    vl_logic;
        PCL_wbClearTerms: out    vl_logic;
        dcdMultiple     : out    vl_logic;
        dcdStringIndexed: out    vl_logic;
        PCL_dIcmpForStuff: out    vl_logic;
        IFB_stuffStL2   : in     vl_logic;
        PCL_sdqMuxSel   : out    vl_logic;
        PCL_wbStrgEnd   : in     vl_logic;
        DBG_exeIacSuppress: in     vl_logic;
        plaMrSel        : in     vl_logic;
        plaMdSel        : in     vl_logic;
        PCL_dcdMrSelQ   : out    vl_logic;
        PCL_dcdMdSelQ   : out    vl_logic;
        PCL_mmuExeAbort : out    vl_logic;
        PCL_wbAlgnErr   : in     vl_logic;
        DBG_wbDacSuppress: in     vl_logic;
        VCT_exeSuppForApu: in     vl_logic;
        exeMmuOp        : in     vl_logic;
        PCL_exeLoadUseHold: out    vl_logic;
        PCL_holdMdMr    : out    vl_logic;
        PCL_exeSrmBpSel : in     vl_logic_vector(0 to 2);
        plaStwcx        : in     vl_logic;
        exeLwarx        : in     vl_logic;
        PCL_dIcmpForWbFlushQDlydL2: out    vl_logic;
        exeRpEqexe2RpAddr: in     vl_logic;
        exeMorMRpEqwbLpAddr: in     vl_logic;
        exeMorMRpEqlwbLpAddr: in     vl_logic;
        VCT_exeSuppForExe2Clear: in     vl_logic;
        wbByteEn        : in     vl_logic_vector(0 to 3);
        DCU_carByteEn   : in     vl_logic_vector(0 to 3);
        PCL_dvcByteEnL2 : out    vl_logic_vector(0 to 3);
        PCL_aRegForEaE2 : out    vl_logic;
        PCL_bRegForEaE2 : out    vl_logic;
        PCL_apuWbHold   : out    vl_logic;
        exeApuExeWbLdUseL2: in     vl_logic;
        exeApuExeLwbLdUseL2: in     vl_logic;
        ltchDA          : out    vl_logic;
        dcdTimSprDcd    : out    vl_logic_vector(0 to 5);
        dcdIcuSprDcd    : out    vl_logic_vector(0 to 2);
        plaMfspr        : in     vl_logic;
        VCT_exeSuppForCr: in     vl_logic;
        dcdDbgSprDcd    : out    vl_logic_vector(0 to 3);
        dcdExeSprDcd    : out    vl_logic_vector(0 to 4);
        dcdVctSprDcd    : out    vl_logic_vector(0 to 5);
        resetL2         : out    vl_logic;
        PCL_dcdLitCntl  : in     vl_logic_vector(2 to 4);
        plaEaCalc       : in     vl_logic;
        exeFullForE1_NEG: in     vl_logic;
        exe2FullForE1_NEG: in     vl_logic;
        wbFullForPO     : in     vl_logic;
        plaApuDiv       : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        PCL_ocmAbortReq : out    vl_logic;
        exeStrgStC0     : in     vl_logic;
        wbLoadForApu    : in     vl_logic;
        PCL_blkFlushForVct: out    vl_logic_vector(0 to 2);
        dcdJtgSprDcd    : out    vl_logic;
        PCL_sraRegE2    : out    vl_logic;
        VCT_sxrOR_L2    : in     vl_logic;
        PCL_exeDvcOrParityHold: out    vl_logic;
        CAR_cacheable   : in     vl_logic;
        PCL_lwbCacheableL2: out    vl_logic;
        PCL_dofDregFull : out    vl_logic;
        ICU_CCR0DPP     : in     vl_logic
    );
end p405s_pipeCntl;
