library verilog;
use verilog.vl_types.all;
entity p405s_apu_shell is
    port(
        clk             : in     vl_logic;
        rst_b           : in     vl_logic;
        C405_apuDcdInstruction: in     vl_logic_vector(0 to 31);
        C405_apuDcdFull : in     vl_logic;
        C405_apuDcdHold : in     vl_logic;
        C405_apuExeHold : in     vl_logic;
        C405_apuExeFlush: in     vl_logic;
        C405_apuExeWdCnt: in     vl_logic_vector(0 to 1);
        C405_apuExeRaData: in     vl_logic_vector(0 to 31);
        C405_apuExeRbData: in     vl_logic_vector(0 to 31);
        C405_apuXerCA   : in     vl_logic;
        C405_apuWbHold  : in     vl_logic;
        C405_apuWbFlush : in     vl_logic;
        C405_apuWbEndian: in     vl_logic;
        C405_apuWbByteEn: in     vl_logic_vector(0 to 3);
        C405_apuExeLoadDBus: in     vl_logic_vector(0 to 31);
        C405_apuExeLoadDValid: in     vl_logic;
        C405_apuMsrFE0  : in     vl_logic;
        C405_apuMsrFE1  : in     vl_logic;
        AltiVec_APU_ValidOp: in     vl_logic;
        AltiVec_APU_ExeBusy: in     vl_logic;
        AltiVec_APU_RaEn: in     vl_logic;
        AltiVec_APU_RbEn: in     vl_logic;
        AltiVec_APU_CR6En: in     vl_logic;
        AltiVec_APU_CRData: in     vl_logic_vector(0 to 3);
        APU_c405DcdValidOp: out    vl_logic;
        APU_c405DcdApuOp: out    vl_logic;
        APU_c405DcdFpuOp: out    vl_logic;
        APU_c405DcdPrivOp: out    vl_logic;
        APU_c405DcdGprWrite: out    vl_logic;
        APU_c405DcdRaEn : out    vl_logic;
        APU_c405DcdRbEn : out    vl_logic;
        APU_c405DcdXerOVEn: out    vl_logic;
        APU_c405DcdXerCAEn: out    vl_logic;
        APU_c405DcdCREn : out    vl_logic;
        APU_c405ExeCRField: out    vl_logic_vector(0 to 2);
        APU_c405DcdForceAlgn: out    vl_logic;
        APU_c405DcdLoad : out    vl_logic;
        APU_c405DcdStore: out    vl_logic;
        APU_c405DcdUpdate: out    vl_logic;
        APU_c405DcdLdStByte: out    vl_logic;
        APU_c405DcdLdStHw: out    vl_logic;
        APU_c405DcdLdStWd: out    vl_logic;
        APU_c405DcdLdStDw: out    vl_logic;
        APU_c405DcdLdStQw: out    vl_logic;
        APU_c405DcdTrapBE: out    vl_logic;
        APU_c405DcdTrapLE: out    vl_logic;
        APU_c405DcdForceBESteering: out    vl_logic;
        APU_c405ExeLdDepend: out    vl_logic;
        APU_c405WbLdDepend: out    vl_logic;
        APU_c405LwbLdDepend: out    vl_logic;
        APU_c405ExeBlockingMCO: out    vl_logic;
        APU_c405ExeNonBlockingMCO: out    vl_logic;
        APU_c405ExeBusy : out    vl_logic;
        APU_c405ExeResult: out    vl_logic_vector(0 to 31);
        APU_c405ExeXerCA: out    vl_logic;
        APU_c405ExeXerOV: out    vl_logic;
        APU_c405ExeCR   : out    vl_logic_vector(0 to 3);
        APU_c405Exception: out    vl_logic;
        APU_c405FpuException: out    vl_logic;
        APU_c405SleepReq: out    vl_logic;
        APU_AltiVec_Ins : out    vl_logic_vector(0 to 31);
        APU_AltiVec_RaData: out    vl_logic_vector(0 to 31);
        APU_AltiVec_RbData: out    vl_logic_vector(0 to 31);
        APU_AltiVec_DcdHold: out    vl_logic
    );
end p405s_apu_shell;
