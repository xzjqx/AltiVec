library verilog;
use verilog.vl_types.all;
entity p405s_storage is
    port(
        PCL_addFour     : out    vl_logic;
        PCL_apuExeWdCnt : out    vl_logic_vector(0 to 1);
        PCL_dcuByteEn   : out    vl_logic_vector(0 to 3);
        PCL_dsOcmByteEn : out    vl_logic_vector(0 to 3);
        PCL_exeEaQwEn   : out    vl_logic_vector(0 to 3);
        algnErr         : out    vl_logic;
        blkExeSpAddr    : out    vl_logic;
        byteCount       : out    vl_logic_vector(6 to 7);
        cntGtEq4        : out    vl_logic;
        exeStrgSt       : out    vl_logic_vector(0 to 2);
        exeStrgStC0     : out    vl_logic;
        sPortSelInc     : out    vl_logic;
        strgEnd         : out    vl_logic;
        strgLpWrEn      : out    vl_logic;
        APU_dcdLdStByte : in     vl_logic;
        APU_dcdLdStDw   : in     vl_logic;
        APU_dcdLdStHw   : in     vl_logic;
        APU_dcdLdStQw   : in     vl_logic;
        APU_dcdLdStWd   : in     vl_logic;
        CB              : in     vl_logic;
        EXE_ea          : in     vl_logic_vector(30 to 31);
        EXE_xerTBC      : in     vl_logic_vector(0 to 6);
        EXE_xerTBCIn    : in     vl_logic_vector(0 to 6);
        IFB_exeFlush    : in     vl_logic;
        PCL_Rbit        : in     vl_logic;
        countE1         : in     vl_logic;
        countE2         : in     vl_logic;
        dcdMultiple     : in     vl_logic;
        dcdRBL2         : in     vl_logic_vector(0 to 4);
        dcdRSRTL2       : in     vl_logic_vector(0 to 4);
        dcdStringImmediate: in     vl_logic;
        dcdStringIndexed: in     vl_logic;
        exeAlg          : in     vl_logic;
        exeApuFpuOp     : in     vl_logic;
        exeByteRev      : in     vl_logic;
        exeDcread       : in     vl_logic;
        exeEaCalc       : in     vl_logic;
        exeForceAlgn    : in     vl_logic;
        exeLd           : in     vl_logic;
        exeLwarx        : in     vl_logic;
        exeMultiple     : in     vl_logic;
        exeStore        : in     vl_logic;
        exeString       : in     vl_logic;
        exeStwcx        : in     vl_logic;
        exeXerTBCUpdInstr: in     vl_logic;
        gtErr           : in     vl_logic;
        nopStringIndexed: in     vl_logic;
        plaApuLdSt      : in     vl_logic;
        plaLdStByte     : in     vl_logic;
        plaLdStDw       : in     vl_logic;
        plaLdStHw       : in     vl_logic;
        plaLdStQw       : in     vl_logic;
        plaLdStWd       : in     vl_logic;
        plaVal          : in     vl_logic;
        storageStMachE1 : in     vl_logic;
        storageStMachE2 : in     vl_logic
    );
end p405s_storage;
