library verilog;
use verilog.vl_types.all;
entity p405s_trcCntlEqs is
    port(
        TRC_se          : out    vl_logic;
        TRC_sleepReq    : out    vl_logic;
        TRC_fifoOneEntryFree: out    vl_logic;
        trcSECtrReset   : out    vl_logic;
        trcReset        : out    vl_logic;
        nxtFifoWrAddr   : out    vl_logic_vector(0 to 3);
        nxtFifoRdAddr   : out    vl_logic_vector(0 to 3);
        nxtFifoStatus   : out    vl_logic_vector(0 to 4);
        nxtTrcSerState  : out    vl_logic_vector(0 to 3);
        nxtTSBus        : out    vl_logic_vector(0 to 3);
        nxtOddCycle     : out    vl_logic;
        nxtStampInc     : out    vl_logic;
        nxtSeCtrEqZero  : out    vl_logic;
        trcESTSE1       : out    vl_logic;
        trcTimeStampE1  : out    vl_logic;
        trcSECtrE1      : out    vl_logic;
        fifoCntlE2      : out    vl_logic;
        serializerE1    : out    vl_logic;
        trcTimeStampE2  : out    vl_logic;
        evenESTEE1      : out    vl_logic;
        trcFifoE1       : out    vl_logic_vector(0 to 15);
        xxxTEQ          : out    vl_logic;
        ICU_traceEnable : in     vl_logic;
        IFB_postEntry   : in     vl_logic;
        IFB_stopAck     : in     vl_logic;
        IFB_seIdleSt    : in     vl_logic;
        VCT_msrWE       : in     vl_logic;
        JTG_stopReq     : in     vl_logic;
        DBG_stopReq     : in     vl_logic;
        XXX_TE          : in     vl_logic;
        serDataOut      : in     vl_logic_vector(0 to 2);
        seInc           : in     vl_logic_vector(0 to 10);
        trcFifoDataOut  : in     vl_logic_vector(30 to 31);
        fifoStatusL2    : in     vl_logic_vector(0 to 4);
        fifoWrAddrL2    : in     vl_logic_vector(0 to 3);
        fifoRdAddrL2    : in     vl_logic_vector(0 to 3);
        trcSerStateL2   : in     vl_logic_vector(0 to 3);
        coreResetL2     : in     vl_logic;
        evenTEL2        : in     vl_logic;
        stampIncL2      : in     vl_logic;
        trcEnableDlyL2  : in     vl_logic;
        oddCycleL2      : in     vl_logic;
        seCtrEqZeroL2   : in     vl_logic;
        xxxTraceDisableL2: in     vl_logic
    );
end p405s_trcCntlEqs;
