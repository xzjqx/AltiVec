// 
// ************************************************************************** 
// 
//  Copyright (c) International Business Machines Corporation, 2005. 
// 
//  This file contains trade secrets and other proprietary and confidential 
//  information of International Business Machines Corporation which are 
//  protected by copyright and other intellectual property rights and shall 
//  not be reproduced, transferred to other documents, disclosed to others, 
//  or used for any purpose except as specifically authorized in writing by 
//  International Business Machines Corporation. This notice must be 
//  contained as part of this text at all times. 
// 
// ************************************************************************** 
//
module p405s_cpu_top( C405_jtgCaptureDR, C405_jtgExtest, C405_jtgPlbDcuPriorityAdjust,
     C405_jtgShiftDR, C405_jtgTDO, C405_jtgTDOEn, C405_jtgUpdateDR, C405_rstChipResetReq,
     C405_rstCoreResetReq, C405_rstSystemResetReq, CPU_TEType, Core_lssdScanOut,
     DCU_parityError, DCU_FlushParityError, EXE_apuLoadData, EXE_dcrAddr, EXE_dcrDataBus, EXE_dcuData,
     EXE_dsEA_NEG, EXE_dsEaCP, EXE_eaARegBuf, EXE_eaBRegBuf,
     EXE_icuSprDcds, EXE_mmuIcuSprDataBus, EXE_raData, EXE_rbData,
     ICU_parityErrE, ICU_parityErrO, ICU_tagParityErr, ICU_CCR0DPP, ICU_CCR0DPE, ICU_CCR0IPE, ICU_CCR0TPE,
     EXE_sprAddr, EXE_xerCa, IFB_TE, IFB_cntxSync, IFB_cntxSyncOCM, IFB_coreSleepReq,
     IFB_dcdFullApuL2, IFB_exeFlush, IFB_extStopAck, IFB_fetchReq, IFB_icuCancelDataL2,
     IFB_isAbortForICU, IFB_isAbortForMMU, IFB_isEA, IFB_isNL, IFB_isNP,
     IFB_isOcmAbus_Neg, IFB_nonSpecAcc, IFB_ocmAbort, IFB_regDcdApuL2,
     IFB_wbIar, JTG_iCacheWr, JTG_instBuf, MMU_tlbREParityErr, MMU_tlbSXParityErr,
     MMU_dsParityErr, MMU_isParityErr, PCL_apuExeWdCnt, PCL_apuLoadDV,
     PCL_apuWbHold, PCL_dcdHoldForApu, PCL_dcuByteEn, PCL_dcuOp,
     PCL_dcuOp_early, PCL_dsMmuOp, PCL_dsOcmByteEn, PCL_exeAbort,
     PCL_exeFlushForApu, PCL_exeHoldForApu, PCL_exeLdNotSt, PCL_exeStorageOp,
     PCL_exeStringMultiple, PCL_exeTlbOp, PCL_icuOp, PCL_mfDCR, PCL_mfSPR,
     PCL_mmuExeAbort, PCL_mmuIcuSprHold, PCL_mmuSprDcd, PCL_mtDCR, PCL_mtSPR,
     PCL_ocmAbortReq, PCL_stSteerCntl, PCL_tlbRE, PCL_tlbSX, PCL_tlbWE, PCL_tlbWS,
     PCL_trcLoadDV, PCL_wbComplete, PCL_wbFull, PCL_wbHoldNonErr, PCL_wbStorageOp,
     TIM_timerResetL2, TRC_evenESBusL2, TRC_oddCycle, TRC_oddESBusL2,
     TRC_tsBusL2, VCT_apuWbFlush, VCT_dcuWbAbort, VCT_dearE2, VCT_errorOut,
     VCT_icuWbAbort, VCT_mmuExeSuppress, VCT_mmuWbAbort, VCT_msrCE, VCT_msrDR, VCT_msrEE,
     VCT_msrFE0, VCT_msrFE1, VCT_msrIR, VCT_msrPR, VCT_msrWE, VCT_timerIntrp, APU_dcdApuOp,
     APU_dcdExeLdDepend, APU_dcdForceAlgn, APU_dcdForceBESteering, APU_dcdFpuOp, APU_dcdGprWr,
     APU_dcdLdStByte, APU_dcdLdStDw, APU_dcdLdStHw, APU_dcdLdStQw, APU_dcdLdStWd, APU_dcdLoad,
     APU_dcdLwbLdDepend, APU_dcdPrivOp, APU_dcdRaEn, APU_dcdRbEn, APU_dcdRc, APU_dcdStore,
     APU_dcdTrapBE, APU_dcdTrapLE, APU_dcdUpdate, APU_dcdValidOp, APU_dcdWbLdDepend,
     APU_dcdXerCAEn, APU_dcdXerOVEn, APU_exception, APU_exeBlkingMco, APU_exeBusy, APU_exeCa,
     APU_exeCr, APU_exeCrField, APU_exeNonBlkingMco, APU_exeOv, APU_exeResult,
     APU_sleepReq, C405_timerTick, CAR_cacheable, CAR_endian, CB, TimerClk, CPM_coreClkOff, DBG_c405DebugHalt,
     DBG_c405ExtBusHoldAck, DCU_CA, DCU_DA, DCU_SCL2, DCU_SDQ_mod, DCU_carByteEn,
     DCU_data_NEG, DCU_diagBus, DCU_firstCycCarStXltV, DCU_pclOcmWait,
     DCU_sleepReq, EIC_critIntrp, EIC_extIntrp, FPU_exception, ICU_EO, ICU_GPRC, ICU_LDBE,
     ICU_diagBus, ICU_dsCA, ICU_ifbError, ICU_isBus, ICU_isCA, ICU_sleepReq,
     ICU_sprDataBus, ICU_syncAfterReset, ICU_traceEnable, JTG_c405BndScanTDO,
     JTG_c405TCK, JTG_c405TDI, JTG_c405TMS, JTG_c405TRST_NEG, 
     LSSD_coreScanIn, LSSD_coreTestEn, LSSD_jtgCClk, MMU_BMCO,
     MMU_dsStateBorC, MMU_dsStatus, MMU_isStatus, MMU_sprDataBus, MMU_tlbSXHit,
     MMU_wbHold, OCM_DOF, OCM_dsComplete, OCM_dsData, PGM_coprocPresent, PGM_dcu_DOF,
     PGM_deterministicMult, PGM_divEn, PGM_mmuEn, PGM_pvrBus, PLB_dcuErr,
     RST_c405ResetChip, RST_c405ResetSystem, TRC_c405TE, TRC_c405TraceDisable, XXX_dcrAck,
     XXX_dcrDataBus, XXX_uncondEvent, c2Clk, resetCore, 
     EXE_gprSysClkPI);
     
output  C405_jtgCaptureDR, C405_jtgExtest, C405_jtgPlbDcuPriorityAdjust, C405_jtgShiftDR,
     C405_jtgTDO, C405_jtgTDOEn, C405_jtgUpdateDR, C405_rstChipResetReq, C405_rstCoreResetReq,
     C405_rstSystemResetReq, EXE_xerCa, IFB_TE, IFB_cntxSync, IFB_cntxSyncOCM,
     IFB_coreSleepReq, IFB_dcdFullApuL2, IFB_exeFlush, IFB_extStopAck, IFB_fetchReq,
     IFB_icuCancelDataL2, IFB_isAbortForMMU, IFB_isNL, IFB_isNP, IFB_nonSpecAcc, IFB_ocmAbort,
     JTG_iCacheWr, PCL_apuLoadDV, PCL_apuWbHold, PCL_dcdHoldForApu, PCL_exeAbort,
     PCL_exeFlushForApu, PCL_exeHoldForApu, PCL_exeLdNotSt, PCL_exeStorageOp,
     PCL_exeStringMultiple, PCL_exeTlbOp, PCL_mfDCR, PCL_mfSPR, PCL_mmuExeAbort,
     PCL_mmuIcuSprHold, PCL_mtDCR, PCL_mtSPR, PCL_ocmAbortReq, PCL_tlbRE, PCL_tlbSX, PCL_tlbWE,
     PCL_tlbWS, PCL_trcLoadDV, PCL_wbComplete, PCL_wbFull, PCL_wbHoldNonErr, PCL_wbStorageOp,
     TIM_timerResetL2, TRC_oddCycle, VCT_apuWbFlush, VCT_dcuWbAbort, VCT_dearE2, VCT_errorOut,
     VCT_icuWbAbort, VCT_mmuExeSuppress, VCT_mmuWbAbort, VCT_msrCE, VCT_msrDR, VCT_msrEE,
     VCT_msrFE0, VCT_msrFE1, VCT_msrIR, VCT_msrPR, VCT_msrWE, VCT_timerIntrp;


input  APU_dcdApuOp, APU_dcdExeLdDepend, APU_dcdForceAlgn, APU_dcdForceBESteering,
     APU_dcdFpuOp, APU_dcdGprWr, APU_dcdLdStByte, APU_dcdLdStDw, APU_dcdLdStHw, APU_dcdLdStQw,
     APU_dcdLdStWd, APU_dcdLoad, APU_dcdLwbLdDepend, APU_dcdPrivOp, APU_dcdRaEn, APU_dcdRbEn,
     APU_dcdRc, APU_dcdStore, APU_dcdTrapBE, APU_dcdTrapLE, APU_dcdUpdate, APU_dcdValidOp,
     APU_dcdWbLdDepend, APU_dcdXerCAEn, APU_dcdXerOVEn, APU_exception, APU_exeBlkingMco,
     APU_exeBusy, APU_exeCa, APU_exeNonBlkingMco, APU_exeOv, APU_sleepReq, C405_timerTick,
     CAR_cacheable, CAR_endian, CPM_coreClkOff, DBG_c405DebugHalt, DBG_c405ExtBusHoldAck, DCU_CA, DCU_DA,
     DCU_parityError, DCU_FlushParityError, DCU_SCL2, DCU_firstCycCarStXltV, DCU_pclOcmWait, DCU_sleepReq, EIC_critIntrp,
     ICU_parityErrE, ICU_parityErrO, ICU_tagParityErr, ICU_CCR0DPP, ICU_CCR0DPE, ICU_CCR0IPE, ICU_CCR0TPE,
     EIC_extIntrp, FPU_exception, ICU_GPRC, ICU_LDBE, ICU_dsCA, ICU_isCA, ICU_sleepReq,
     ICU_syncAfterReset, ICU_traceEnable, JTG_c405BndScanTDO, JTG_c405TCK, JTG_c405TDI,
     JTG_c405TMS, JTG_c405TRST_NEG, LSSD_coreTestEn, LSSD_jtgCClk,
     MMU_BMCO, MMU_dsStateBorC, MMU_tlbREParityErr, MMU_tlbSXParityErr,
     MMU_dsParityErr, MMU_isParityErr, MMU_tlbSXHit, MMU_wbHold, OCM_DOF,
     OCM_dsComplete, PGM_coprocPresent, PGM_dcu_DOF, PGM_deterministicMult, PGM_divEn,
     PGM_mmuEn, PLB_dcuErr, RST_c405ResetChip, RST_c405ResetSystem, TRC_c405TE,
     TRC_c405TraceDisable, XXX_dcrAck, XXX_uncondEvent, c2Clk, resetCore;

// added for tbird
input	       EXE_gprSysClkPI;


output [0:31]  EXE_apuLoadData;
output [0:31]  EXE_raData;
output [0:31]  IFB_regDcdApuL2;
output [0:9]  PCL_stSteerCntl;
output [0:1]  TRC_oddESBusL2;
output [0:31]  EXE_dsEA_NEG;
output [0:3]  PCL_dsMmuOp;
output [0:3]  TRC_tsBusL2;
output [0:29]  IFB_wbIar;
output [0:2]  IFB_isAbortForICU;
output [0:31]  EXE_rbData;
output [0:1]  TRC_evenESBusL2;
output [0:7]  EXE_dsEaCP;
output [0:1]  PCL_apuExeWdCnt;
output [0:29]  IFB_isEA;
output [0:2]  EXE_icuSprDcds;
output [0:3]  PCL_dcuByteEn;
output [0:29]  IFB_isOcmAbus_Neg;
output [0:21]  EXE_eaBRegBuf;
output [0:31]  EXE_dcuData;
output [0:2]  PCL_dcuOp_early;
output [0:3]  PCL_dsOcmByteEn;
output [0:11]  PCL_dcuOp;
output [0:21]  EXE_eaARegBuf;
output [0:31]  EXE_dcrDataBus;
output [0:31]  EXE_mmuIcuSprDataBus;
output [4:9]  EXE_sprAddr;
output [0:31]  JTG_instBuf;
output [0:10]  CPU_TEType;
output [0:8]  PCL_mmuSprDcd;
output [0:9]  EXE_dcrAddr;
output [0:3]  PCL_icuOp;
output [10:31]  Core_lssdScanOut;


input [0:1]  MMU_isStatus;
input [0:31]  PGM_pvrBus;
input [0:31]  XXX_dcrDataBus;
input [0:31]  OCM_dsData;
input [0:1]  ICU_ifbError;
input [0:31]  ICU_sprDataBus;
input [0:31]  APU_exeResult;
input [0:31]  MMU_sprDataBus;
input [0:3]  DCU_carByteEn;
input [0:31]  DCU_data_NEG;
input [0:31]  DCU_SDQ_mod;
input [0:2]  APU_exeCrField;
input [0:3]  APU_exeCr;
input [0:22]  ICU_diagBus;
input [0:63]  ICU_isBus;
input [0:1]  ICU_EO;
input [0:20]  DCU_diagBus;
input CB;
input TimerClk;
input [0:7]  MMU_dsStatus;
input [10:31]  LSSD_coreScanIn;

// Buses in the design
wire  [0:3]  PCL_exeRbEn;
wire  [0:31] EXE_vctDbgSprDataBus;
wire  [0:3]  PCL_dvcByteEnL2;
wire  [0:2]  DBG_immdTE;
wire  [0:31] JTG_sprDataBus;
wire  [0:7]  VCT_vectorBus;
wire  [0:31] VCT_sprDataBus;
wire  [0:31] DBG_sprDataBus;
wire  [0:2]  PCL_dcdHoldForIfb;
wire  [0:4]  PCL_exeTrapCond;
wire  [0:3]  EXE_cc;
wire  [0:6]  EXE_xerTBCIn;
wire  [0:31] IFB_dcdDataIn_Neg;
wire  [0:7]  PCL_ldMuxSel;
wire  [0:9]  PCL_dcdSpAddr;
wire  [0:4]  PCL_wbRpAddr;
wire  [0:7]  PCL_ldSteerMuxSel;
wire  [0:1]  PCL_exe2AccRegMuxSel;
wire  [0:2]  PCL_blkFlushForVct;
wire  [0:29] IFB_traceData;
wire  [0:31] JTG_inst;
wire  [30:31]EXE_ea;
wire  [0:9]  PCL_dcdApAddr;
wire  [0:31] TIM_sprDataBus;
wire  [0:3]  EXE_dvc2ByteCmp;
wire  [0:3]  PCL_exeAdmCntl;
wire  [0:1]  PCL_ldAdjMuxSel;
wire  [0:1]  PCL_exe2MacOrMultEnForMS;
wire  [0:31] EXE_ifbSprDataBus;
wire  [0:4]  DBG_wbTE;
wire  [0:1]  PCL_exeMultEn_NEG;
wire  [0:4]  PCL_exeSprDcds;
wire  [0:3]  PCL_dbgSprDcds;
wire  [0:5]  PCL_timSprDcds;
wire  [0:2]  PCL_srmRegE2;
wire  [0:31] EXE_timJtgSprDataBus;
wire  [0:3]  PCL_exeSrmCntl;
wire  [0:2]  EXE_xer;
wire  [0:1]  EXE_gprSO;
wire  [0:3]  PCL_exeRaEn;
wire  [0:4]  DBG_exeTE;
wire  [0:9]  PCL_dcdBpAddr;
wire  [0:1]  IFB_dcdFullL2;
wire  [0:4]  PCL_dcdLitCntl;
wire  [0:4]  PCL_lwbLpAddr;
wire  [0:6]  EXE_xerTBC;
wire  [0:2]  PCL_exeSrmBpSel;
wire  [0:1]  PCL_exeDivEnForMuxSel;
wire  [1:3]  PCL_ldAdjG1;
wire  [0:4]  IFB_exeIfetchErrL2;
wire  [0:9]  PCL_diagBus;
wire  [0:5]  PCL_vctSprDcds;
wire  [0:3]  EXE_dvc1ByteCmp;
wire  [11:31]PCL_dcdImmd;
wire  [0:5]  PCL_ldFillByPassMuxSel;
wire  [0:3]  PCL_exeEaQwEn;
wire  [0:2]  PCL_dcdSrmMuxSel;
wire  [0:11] VCT_sxr;
wire  [0:31] IFB_sprDataBus;
wire  [0:1]  PCL_dofDregMuxSel;
wire  [0:7]  PCL_exeLogicalCntl;
wire  [0:1]  PCL_exeMultEnForMuxSel;
wire  [0:1]  PCL_exeAddSgndOp_NEG;
wire  [0:1]  IFB_traceType;
wire  [0:1]  PCL_exe2MacOrMultEn_NEG;
wire  [1:2]  IFB_traceESL2;
wire  [0:7]  IFB_diagBus;

wire         PCL_gprRdClk;
wire dcdApuValidOp_NEG;


// Replacing instantiation: INVERT I1428
assign dcdApuValidOp_NEG = ~(APU_dcdValidOp);


p405s_jtg_top
 jtg_topSch(
        .JTG_TDO(                           C405_jtgTDO),
        .JTG_captureDR(                     C405_jtgCaptureDR),
        .JTG_dbdrPulse(                     JTG_dbdrPulse),
        .JTG_dbgWaitEn(                     JTG_dbgWaitEn),
        .JTG_extest(                        C405_jtgExtest),
        .JTG_freezeTimers(                  JTG_freezeTimers),
        .JTG_iCacheWr_NEG(                  JTG_iCacheWr),
        .JTG_inst(                          JTG_inst[0:31]),
        .JTG_instBuf(                       JTG_instBuf[0:31]),
        .JTG_pgmOut(                        C405_jtgPlbDcuPriorityAdjust),
        .JTG_resetChipReq(                  C405_rstChipResetReq),
        .JTG_resetCoreReq(                  C405_rstCoreResetReq),
        .JTG_resetDBSR(                     JTG_resetDbsr),
        .JTG_resetSystemReq(                C405_rstSystemResetReq),
        .JTG_shiftDR(                       C405_jtgShiftDR),
        .JTG_sprDataBus(                    JTG_sprDataBus[0:31]),
        .JTG_step(                          JTG_step),
        .JTG_stepUPD(                       JTG_stepUPD),
        .JTG_stopReq(                       JTG_stopReq),
        .JTG_stuff(                         JTG_stuff),
        .JTG_stuffUPD(                      JTG_stuffUPD),
        .JTG_tDOEnable(                     C405_jtgTDOEn),
        .JTG_uncondEvent(                   JTG_uncondEvent),
        .JTG_updateDR(                      C405_jtgUpdateDR),
        .CB(                                CB),
        .CPM_coreClkOff(                    CPM_coreClkOff),
        .DBG_DE(                            DBG_eventSet),
        .DBG_UDE(                           DBG_udeEventSet),
        .DBG_resetChip(                     DBG_resetChip),
        .DBG_resetCore(                     DBG_resetCore),
        .DBG_resetSystem(                   DBG_resetSystem),
        .EXE_sprDataBus(                    EXE_timJtgSprDataBus[0:31]),
        .ICU_sleepReq(                      ICU_sleepReq),
        .IFB_msrWE(                         VCT_msrWEL2),
        .IFB_rstStepPend(                   IFB_rstStepPend),
        .IFB_rstStuffPend(                  IFB_rstStuffPend),
        .IFB_stopAck(                       IFB_stopAck),
        .JTGEX_BndScanTDO(                  JTG_c405BndScanTDO),
        .JTGEX_TCK(                         JTG_c405TCK),
        .JTGEX_TDI(                         JTG_c405TDI),
        .JTGEX_TMS(                         JTG_c405TMS),
        .JTGEX_TRST_NEG(                    JTG_c405TRST_NEG),
        .PCL_exeMfspr(                      PCL_mfSPR),
        .PCL_exeMtspr(                      PCL_mtSPR),
        .PCL_exeSprHold(                    PCL_timJtgsprHold),
        .PCL_jtgSprDcd(                     PCL_jtgSprDcd),
        .PLB_jtgHoldAck(                    DBG_c405ExtBusHoldAck),
        .TIM_wdChipRst(                     TIM_wdChipRst),
        .TIM_wdCoreRst(                     TIM_wdCoreRst),
        .TIM_wdSysRst(                      TIM_wdSysRst),
        .VCT_msrDWE(                        VCT_msrDWE),
        .VCT_srr1DWE(                       VCT_srr1DWE),
        .VCT_srr3DWE(                       VCT_srr3DWE),
        .VCT_stuffStepSup(                  VCT_stuffStepSup),
        .VCT_sxr(                           VCT_sxr[0:11]),
        .XXX_coreReset(                     resetCore),
        .XXX_jtgHalt(                       DBG_c405DebugHalt),
        .XXX_systemReset(                   RST_c405ResetSystem),
        .jtgDiagBus1(                       {PCL_diagBus[0:9], IFB_diagBus[0:7], 1'b0,
                                             1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
                                             1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
                                             1'b0, 1'b0, 1'b0}),
        .jtgDiagBus2(                       {ICU_diagBus[0:22],
                                             1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
                                             1'b0, 1'b0, 1'b0, 1'b0}),
        .jtgDiagBus3(                       {DCU_diagBus[0:20], 1'b0, 1'b0, 1'b0,
                                             1'b0, 1'b0, 1'b0, 1'b0,
                                             1'b0, 1'b0, 1'b0, 1'b0})
         );

p405s_dbg_top
 dbg_topSch(
        .DBG_dacEn(                         DBG_dacEn),
        .DBG_dacIntrp(                      symNet480),
        .DBG_dvcRdEn(                       DBG_dvcRdEn),
        .DBG_dvcWrEn(                       DBG_dvcWrEn),
        .DBG_eventSet(                      DBG_eventSet),
        .DBG_exeIacSuppress(                DBG_exeIacSuppress),
        .DBG_exeSuppress(                   DBG_exeSuppress),
        .DBG_exeTE(                         DBG_exeTE[0:4]),
        .DBG_freezeTimers(                  DBG_freezeTimers),
        .DBG_iacEn(                         DBG_iacEn),
        .DBG_icmpEn(                        DBG_icmpEn),
        .DBG_immdTE(                        DBG_immdTE[0:2]),
        .DBG_intrp(                         DBG_intrp),
        .DBG_rstChipReq(                    DBG_resetChip),
        .DBG_rstCoreReq(                    DBG_resetCore),
        .DBG_rstSystemReq(                  DBG_resetSystem),
        .DBG_sprDataBus(                    DBG_sprDataBus[0:31]),
        .DBG_stopReq(                       DBG_stopReq),
        .DBG_trapEnQ(                       DBG_trapEnQ),
        .DBG_udeEventSet(                   DBG_udeEventSet),
        .DBG_udeIntrp(                      DBG_udeIntrp),
        .DBG_wbDacSuppress(                 DBG_wbDacSuppress),
        .DBG_wbTE(                          DBG_wbTE[0:4]),
        .DBG_weakStopReq(                   DBG_weakStopReq),
        .CB(                                CB),
        .EXE_dac1Bits0to26Eq(               EXE_dac1Bits0to26Eq),
        .EXE_dac1Bits27to29Eq(              EXE_dac1Bits27to29Eq),
        .EXE_dac1Bits30Eq(                  EXE_dac1Bits30Eq),
        .EXE_dac1Bits31Eq(                  EXE_dac1Bits31Eq),
        .EXE_dac1GtDsEa(                    EXE_dac1GtDsEa),
        .EXE_dac2Bits0to26Eq(               EXE_dac2Bits0to26Eq),
        .EXE_dac2Bits27to29Eq(              EXE_dac2Bits27to29Eq),
        .EXE_dac2Bits30Eq(                  EXE_dac2Bits30Eq),
        .EXE_dac2Bits31Eq(                  EXE_dac2Bits31Eq),
        .EXE_dac2GtDsEa(                    EXE_dac2GtDsEa),
        .EXE_dbgSprDcds(                    PCL_dbgSprDcds[0:3]),
        .EXE_dvc1ByteCmp(                   EXE_dvc1ByteCmp[0:3]),
        .EXE_dvc2ByteCmp(                   EXE_dvc2ByteCmp[0:3]),
        .EXE_sprDataBus(                    EXE_vctDbgSprDataBus[0:31]),
        .IFB_dcdFullL2(                     IFB_dcdFullL2[1]),
        .IFB_exeBrTaken(                    IFB_dbgBrTaken),
        .IFB_exeClear(                      IFB_exeClear),
        .IFB_exeDisableDbL2(                IFB_exeDisalbeDbL2),
        .IFB_exeFlush(                      IFB_exeFlush),
        .IFB_exeFullL2(                     IFB_exeFullL2),
        .IFB_iac1BitsEq(                    IFB_iac1BitsEq),
        .IFB_iac1GtIar(                     IFB_iac1GtIar),
        .IFB_iac2BitsEq(                    IFB_iac2BitsEq),
        .IFB_iac2GtIar(                     IFB_iac2GtIar),
        .IFB_iac3BitsEq(                    IFB_iac3BitsEq),
        .IFB_iac3GtIar(                     IFB_iac3GtIar),
        .IFB_iac4BitsEq(                    IFB_iac4BitsEq),
        .IFB_iac4GtIar(                     IFB_iac4GtIar),
        .IFB_stuffStL2(                     IFB_stuffStL2),
        .IFB_wbDisableDbL2(                 IFB_wbDisalbeDbL2),
        .JTG_dbdrPulse(                     JTG_dbdrPulse),
        .JTG_dbgWaitEn(                     JTG_dbgWaitEn),
        .JTG_resetDBSR(                     JTG_resetDbsr),
        .JTG_uncondEvent(                   JTG_uncondEvent),
        .PCL_dvcCmpEn(                      PCL_dvcCmpEn),
        .PCL_exeDbgLdOp(                    PCL_exeDbgLdOp),
        .PCL_exeDbgRdOp(                    PCL_exeDbgRdOp),
        .PCL_exeDbgStOp(                    PCL_exeDbgStOp),
        .PCL_exeDbgWrOp(                    PCL_exeDbgWrOp),
        .PCL_exeDvcHold(                    PCL_exeDvcHold),
        .PCL_exeIarHold(                    PCL_exeIarHold),
        .PCL_exeTrap(                       PCL_exeTrap),
        .PCL_mtSPR(                         PCL_mtSPR),
        .PCL_sprHold(                       PCL_vctDbgsprHold),
        .PCL_wbClearOrFlush(                PCL_wbClear),
        .PCL_wbDbgIcmp(                     PCL_wbDbgIcmp),
        .PCL_wbFull(                        PCL_wbFullL2),
        .PCL_wbHold(                        PCL_wbHold),
        .VCT_exeBrTrapErrSuppress(          VCT_exeBrTrapErrSuppress),
        .VCT_msrDE(                         VCT_msrDE),
        .VCT_msrDWE(                        VCT_msrDWE),
        .VCT_swapQ01(                       VCT_swapQ01),
        .VCT_swapQ23(                       VCT_swapQ23),
        .VCT_wbErrSuppress(                 VCT_wbErrSuppress),
        .VCT_wbFlush(                       VCT_wbFlush),
        .XXX_uncondEvent(                   XXX_uncondEvent),
        .chipReset(                         RST_c405ResetChip),
        .coreReset(                         resetCore),
        .systemReset(                       RST_c405ResetSystem),
        .PCL_exeDvcOrParityHold(            PCL_exeDvcOrParityHold)            
        );

p405s_trc_top
 trc_topSch(
        .TRC_evenESBusL2(                   TRC_evenESBusL2[0:1]),
        .TRC_fifoFull(                      TRC_fifoFull),
        .TRC_fifoOneEntryFree(              TRC_fifoOneEntryFree),
        .TRC_oddCycleL2(                    TRC_oddCycle),
        .TRC_oddESBusL2(                    TRC_oddESBusL2[0:1]),
        .TRC_se(                            TRC_se),
        .TRC_seCtrEqZeroL2(                 TRC_seCtrEqZeroL2),
        .TRC_sleepReq(                      TRC_sleepReq),
        .TRC_tsBusL2(                       TRC_tsBusL2[0:3]),
        .CB(                                CB),
        .DBG_stopReq(                       DBG_stopReq),
        .ICU_traceEnable(                   ICU_traceEnable),
        .IFB_postEntry(                     IFB_postEntry),
        .IFB_seIdleSt(                      IFB_seIdleSt),
        .IFB_stopAck(                       IFB_stopAck),
        .IFB_traceData(                     IFB_traceData[0:29]),
        .IFB_traceESL2(                     IFB_traceESL2[1:2]),
        .IFB_traceType(                     IFB_traceType[0:1]),
        .JTG_stopReq(                       JTG_stopReq),
        .VCT_msrWE(                         VCT_msrWEL2),
        .XXX_TE(                            TRC_c405TE),
        .XXX_traceDisable(                  TRC_c405TraceDisable),
        .coreReset(                         resetCore)
        );

p405s_vct_top
 vct_topSch(
        .VCT_errorOut(                      VCT_errorOut),
        .VCT_msrDR(                         VCT_msrDR),
        .VCT_msrIR(                         VCT_msrIR),
        .VCT_wbRfci(                        VCT_wbRfci),
        .VCT_wbRfi(                         VCT_wbRfi),
        .VCT_sxr(                           VCT_sxr[0:11]),
        .VCT_swap01(                        VCT_swap01),
        .VCT_swap23(                        VCT_swap23),
        .VCT_vectorBus(                     VCT_vectorBus[0:7]),
        .VCT_msrWE(                         VCT_msrWE),
        .VCT_errorSprSuppress(              VCT_errorSprSuppress),
        .VCT_sprDataBus(                    VCT_sprDataBus[0:31]),
        .VCT_msrDE(                         VCT_msrDE),
        .VCT_swapQ01(                       VCT_swapQ01),
        .VCT_swapQ23(                       VCT_swapQ23),
        .PLB_dcuErr(                        PLB_dcuErr),
        .PCL_wbLdNotSt(                     PCL_wbLdNotSt),
        .PCL_mtSPR(                         PCL_mtSPR),
        .PCL_sprHold(                       PCL_vctDbgsprHold),
        .EIC_critIntrp(                     EIC_critIntrp),
        .EIC_extIntrp(                      EIC_extIntrp),
        .PCL_algnErr(                       PCL_algnErr),
        .ICU_CCR0DPE(                       ICU_CCR0DPE),
        .ICU_CCR0DPP(                       ICU_CCR0DPP),
        .ICU_CCR0IPE(                       ICU_CCR0IPE),
        .ICU_CCR0TPE(                       ICU_CCR0TPE),
        .IFB_exeFlush(                      IFB_exeFlush),
        .PCL_dofDregFull(                   PCL_dofDregFull),
        .PCL_exeCpuOp(                      PCL_exeIllegalOpLtch),
        .IFB_exeIfetchErr(                  IFB_exeIfetchErrL2[0:4]),
        .PCL_exeWrExtEn(                    PCL_exeWrExtEn),
        .PCL_exePrivOp(                     PCL_exePrivOp),
        .PCL_exeDvcOrParityHold(            PCL_exeDvcOrParityHold),
        .PCL_lwbCacheableL2(                PCL_lwbCacheableL2),
        .IFB_stuffStL2(                     IFB_stuffStL2),
        .IFB_swapEnable(                    IFB_swapEnable),
        .IFB_exeISideMachChk(               IFB_exeISideMachChk),
        .CB(                                CB),
        .coreReset(                         resetCore),
        .MMU_dsStatus(                      MMU_dsStatus[0:7]),
        .MMU_dsParityErr(                   MMU_dsParityErr),
        .MMU_tlbSXParityErr(                MMU_tlbSXParityErr),
        .MMU_tlbREParityErr(                MMU_tlbREParityErr),
        .EXE_dofDregParityErrL2(            EXE_dofDregParityErrL2),
        .EXE_wrteeIn(                       EXE_wrteeIn),
        .DBG_intrp(                         DBG_intrp),
        .DBG_exeIacSuppress(                DBG_exeIacSuppress),
        .DBG_trapEnQ(                       DBG_trapEnQ),
        .TIM_fitIntrp(                      TIM_fitIntrp),
        .TIM_pitIntrp(                      TIM_pitIntrp),
        .PCL_exeTrap(                       PCL_exeTrap),
        .TIM_watchDogIntrp(                 TIM_watchDogIntrp),
        .PGM_pvrBus(                        PGM_pvrBus[0:31]),
        .VCT_exeSuppress(                   VCT_exeSuppress),
        .VCT_anySwap(                       VCT_anySwap),
        .PCL_exeApuOp(                      PCL_exeApuOp),
        .DBG_exeSuppress(                   DBG_exeSuppress),
        .VCT_msrCE(                         VCT_msrCE),
        .VCT_msrEE(                         VCT_msrEE),
        .DBG_wbDacSuppress(                 DBG_wbDacSuppress),
        .PCL_exeApuValidOp(                 PCL_exeValidOp),
        .VCT_timerIntrp(                    VCT_timerIntrp),
        .VCT_sxrOR_L2(                      VCTsxrOR_L2),
        .PCL_exeFull(                       PCL_exeFull),
        .JTG_stopReq(                       JTG_stopReq),
        .DBG_stopReq(                       DBG_stopReq),
        .IFB_runStL2(                       IFB_runStL2),
        .APU_exception(                     APU_exception),
        .VCT_msrPR(                         VCT_msrPR),
        .PGM_mmuEn(                         PGM_mmuEn),
        .PCL_dIcmpForWbFlushQDlydL2(        PCL_dIcmpForWbFlushQDlydL2),
        .EXE_vctSprDcds(                    PCL_vctSprDcds[0:5]),
        .EXE_sprDataBus(                    EXE_vctDbgSprDataBus[0:31]),
        .VCT_dcuWbAbort(                    VCT_dcuWbAbort),
        .VCT_wbSuppress(                    VCT_wbSuppress),
        .IFB_exeRfi(                        IFB_exeRfiL2),
        .IFB_exeRfci(                       IFB_exeRfciL2),
        .IFB_exeSc(                         IFB_exeScL2),
        .PCL_wbFull(                        PCL_wbFullL2),
        .VCT_dearE2(                        VCT_dearE2),
        .VCT_wbFlush(                       VCT_wbFlush),
        .PCL_blkFlush(                      PCL_blkFlushForVct[0:2]),
        .VCT_icuWbAbort(                    VCT_icuWbAbort),
        .PCL_exeDvcHold(                    PCL_exeDvcHold),
        .MMU_dsStateBorC(                   MMU_dsStateBorC),
        .PCL_exeFpuOp(                      PCL_exeFpuOp),
        .FPU_exception(                     FPU_exception),
        .PCL_wbHold(                        PCL_wbHold),
        .DBG_udeIntrp(                      DBG_udeIntrp),
        .DBG_weakStopReq(                   DBG_weakStopReq),
        .VCT_msrFE0(                        VCT_msrFE0),
        .VCT_msrFE1(                        VCT_msrFE1),
        .VCT_msrDWE(                        VCT_msrDWE),
        .VCT_wbErrSuppress(                 VCT_wbErrSuppress),
        .VCT_stuffStepSupL2(                VCT_stuffStepSup),
        .VCT_srr1DWE(                       VCT_srr1DWE),
        .VCT_srr3DWE(                       VCT_srr3DWE),
        .IFB_stepStL2(                      IFB_stepStL2),
        .VCT_exeBrTrapErrSuppress(          VCT_exeBrTrapErrSuppress),
        .VCT_wbFlushAsync(                  VCT_wbFlushAsync),
        .VCT_msrWEL2(                       VCT_msrWEL2),
        .PCL_wbStorageOp(                   PCL_wbStorageOp),
        .VCT_wbLoadSuppress(                VCT_wbLoadSuppress),
        .IFB_swapStL2(                      IFB_swapStL2),
        .PCL_exe2Full(                      PCL_exe2Full),
        .JTG_dbgWaitEn(                     JTG_dbgWaitEn),
        .IFB_dcdFullL2(                     IFB_dcdFullL2[1]),
        .VCT_mmuWbAbort(                    VCT_mmuWbAbort),
        .MMU_wbHold(                        MMU_wbHold),
        .VCT_mmuExeSuppress(                VCT_mmuExeSuppress),
        .VCT_exeSuppForApu(                 VCT_exeSuppForApu),
        .DCU_SCL2(                          DCU_SCL2),
        .DCU_FlushParityError(              DCU_FlushParityError),
        .PCL_wbHoldNonErr(                  PCL_wbHoldNonErr),
        .VCT_exeSuppForExe2Clear(           VCT_exeSuppForExe2Clear),
        .VCT_apuWbFlush(                    VCT_apuWbFlush),
        .VCT_exeSuppForCr(                  VCT_exeSuppForCr),
        .LSSD_coreTestEn(                   LSSD_coreTestEn),
        .JTG_stepUPD(                       JTG_stepUPD),
        .JTG_stuffUPD(                      JTG_stuffUPD),
        .lwbFullL2(                         lwbFullL2)
        );

p405s_timer_top
 tim_top(
        .TIM_fitIntrp(                      TIM_fitIntrp),
        .TIM_pitIntrp(                      TIM_pitIntrp),
        .TIM_sprDataBus(                    TIM_sprDataBus[0:31]),
        .TIM_timerResetL2Buf(               TIM_timerResetL2),
        .TIM_watchDogIntrp(                 TIM_watchDogIntrp),
        .TIM_wdChipRst(                     TIM_wdChipRst),
        .TIM_wdCoreRst(                     TIM_wdCoreRst),
        .TIM_wdSysRst(                      TIM_wdSysRst),
        .CB(TimerClk),
        .DBG_freezeTimers(                  DBG_freezeTimers),
        .EXE_sprDataBus(                    EXE_timJtgSprDataBus[0:31]),
        .EXE_timSprDcds(                    PCL_timSprDcds[0:5]),
        .JTG_freezeTimers(                  JTG_freezeTimers),
        .LSSD_coreTestEn(                   LSSD_coreTestEn),
        .OSC_timer(                         C405_timerTick),
        .PCL_mtSPR(                         PCL_mtSPR),
        .PCL_sprHold(                       PCL_timJtgsprHold),
        .resetCore(                         resetCore)
        );

p405s_ifb_top
 ifb_topSch(
        .IFB_TEL2(                          IFB_TE),
        .IFB_TETypeL2(                      CPU_TEType[0:10]),
        .IFB_cntxSync(                      IFB_cntxSync),
        .IFB_cntxSyncOCM(                   IFB_cntxSyncOCM),
        .IFB_coreSleepReqL2(                IFB_coreSleepReq),
        .IFB_dcdApu(                        IFB_regDcdApuL2[0:31]),
        .IFB_dcdBubble(                     IFB_dcdBubble),
        .IFB_dcdDataIn_Neg(                 IFB_dcdDataIn_Neg[0:31]),
        .IFB_dcdFullApuL2(                  IFB_dcdFullApuL2),
        .IFB_dcdFullL2(                     IFB_dcdFullL2[0:1]),
        .IFB_dcdRegE1(                      IFB_dcdRegE1),
        .IFB_dcdRegE2(                      IFB_dcdRegE2),
        .IFB_diagBus(                       IFB_diagBus[0:7]),
        .IFB_exeClear(                      IFB_exeClear),
        .IFB_exeCorrect(                    IFB_exeCorrect),
        .IFB_exeDbgBrTaken(                 IFB_dbgBrTaken),
        .IFB_exeDisableDbL2(                IFB_exeDisalbeDbL2),
        .IFB_exeFlushA(                     IFB_exeFlush),
        .IFB_exeFlushB(                     IFB_exeFlushB),
        .IFB_exeFullL2(                     IFB_exeFullL2),
        .IFB_exeIfetchErrL2(                IFB_exeIfetchErrL2[0:4]),
        .IFB_exeMcrxrL2(                    IFB_exeMcrxrL2),
        .IFB_exeOpForExe2L2(                IFB_exeOpForExe2L2),
        .IFB_exeRfciL2(                     IFB_exeRfciL2),
        .IFB_exeRfiL2(                      IFB_exeRfiL2),
        .IFB_exeScL2(                       IFB_exeScL2),
        .IFB_extStopAck(                    IFB_extStopAck),
        .IFB_fetchReq(                      IFB_fetchReq),
        .IFB_iac1BitsEq(                    IFB_iac1BitsEq),
        .IFB_iac1GtIar(                     IFB_iac1GtIar),
        .IFB_iac2BitsEq(                    IFB_iac2BitsEq),
        .IFB_iac2GtIar(                     IFB_iac2GtIar),
        .IFB_iac3BitsEq(                    IFB_iac3BitsEq),
        .IFB_iac3GtIar(                     IFB_iac3GtIar),
        .IFB_iac4BitsEq(                    IFB_iac4BitsEq),
        .IFB_iac4GtIar(                     IFB_iac4GtIar),
        .IFB_icuCancelDataL2(               IFB_icuCancelDataL2),
        .IFB_isAbortForICU(                 IFB_isAbortForICU[0:2]),
        .IFB_isAbortForMMU(                 IFB_isAbortForMMU),
        .IFB_isEA(                          IFB_isEA[0:29]),
        .IFB_isNL(                          IFB_isNL),
        .IFB_isNP(                          IFB_isNP),
        .IFB_isOcmAbus(                     IFB_isOcmAbus_Neg[0:29]),
        .IFB_nonSpecAcc(                    IFB_nonSpecAcc),
        .IFB_ocmAbort(                      IFB_ocmAbort),
        .IFB_postEntry(                     IFB_postEntry),
        .IFB_rstStepPend(                   IFB_rstStepPend),
        .IFB_rstStuffPend(                  IFB_rstStuffPend),
        .IFB_runStL2(                       IFB_runStL2),
        .IFB_seIdleSt(                      IFB_seIdleSt),
        .IFB_sprDataBus(                    IFB_sprDataBus[0:31]),
        .IFB_stepStL2(                      IFB_stepStL2),
        .IFB_stopAck(                       IFB_stopAck),
        .IFB_stuffStL2(                     IFB_stuffStL2),
        .IFB_swapEnable(                    IFB_swapEnable),
        .IFB_swapStL2(                      IFB_swapStL2),
        .IFB_traceData(                     IFB_traceData[0:29]),
        .IFB_traceESL2(                     IFB_traceESL2[1:2]),
        .IFB_tracePipeHold(                 IFB_tracePipeHold),
        .IFB_traceType(                     IFB_traceType[0:1]),
        .IFB_wbDisableDbL2(                 IFB_wbDisalbeDbL2),
        .IFB_wbIar(                         IFB_wbIar[0:29]),
        .APU_dcdCrField(                    APU_exeCrField[0:2]),
        .APU_dcdRc(                         APU_dcdRc),
        .APU_sleepReq(                      APU_sleepReq),
        .CB(                                CB),
        .DBG_exeTE(                         DBG_exeTE[0:4]),
        .DBG_iacEn(                         DBG_iacEn),
        .DBG_immdTE(                        DBG_immdTE[0:2]),
        .DBG_stopReq(                       DBG_stopReq),
        .DBG_wbTE(                          DBG_wbTE[0:4]),
        .DBG_weakStopReq(                   DBG_weakStopReq),
        .DCU_sleepReq(                      DCU_sleepReq),
        .EXE_cc(                            EXE_cc[0:3]),
        .EXE_sprDataBus(                    EXE_ifbSprDataBus[0:31]),
        .EXE_xer(                           EXE_xer[0:2]),
        .ICU_ifbE(                          ICU_EO[0]),
        .ICU_ifbEDataBus(                   ICU_isBus[0:31]),
        .ICU_ifbError(                      ICU_ifbError[0:1]),
        .ICU_ifbO(                          ICU_EO[1]),
        .ICU_ifbODataBus(                   ICU_isBus[32:63]),
        .ICU_isCA(                          ICU_isCA),
        .ICU_sleepReq(                      ICU_sleepReq),
        .ICU_syncAfterReset(                ICU_syncAfterReset),
        .ICU_traceEnable(                   ICU_traceEnable),
        .JTG_dbdrPulse(                     JTG_dbdrPulse),
        .JTG_inst(                          JTG_inst[0:31]),
        .JTG_step(                          JTG_step),
        .JTG_stopReq(                       JTG_stopReq),
        .JTG_stuff(                         JTG_stuff),
        .LSSD_coreTestEn(                   LSSD_coreTestEn),
        .MMU_isStatus(                      MMU_isStatus[0:1]),
        .MMU_tlbSXHit(                      MMU_tlbSXHit),
        .PCL_Rbit(                          PCL_Rbit),
        .PCL_blkFlush(                      PCL_blkFlush),
        .PCL_dIcmpForStep(                  PCL_dIcmpForStep),
        .PCL_dIcmpForStuff(                 PCL_dIcmpForStuff),
        .PCL_dcdHoldForIFB(                 PCL_dcdHoldForIfb[0:2]),
        .PCL_exe2DataE1(                    PCL_exe2DataE1),
        .PCL_exe2DataE2(                    PCL_exe2DataE2),
        .PCL_exe2FlushorClear(              PCL_exe2FlushorClear),
        .PCL_exe2Full(                      PCL_exe2Full),
        .PCL_exe2IarE1(                     PCL_exe2IarE1),
        .PCL_exe2IarE2(                     PCL_exe2IarE2),
        .PCL_exeHoldForCr(                  PCL_exeHoldForCr),
        .PCL_exeIarHold(                    PCL_exeIarHold),
        .PCL_icuOp_0(                       PCL_icuOp[0]),
        .PCL_sprHold(                       PCL_ifbSprHold),
        .PCL_wbClearTerms(                  PCL_wbClearTerms),
        .PCL_wbFull(                        PCL_wbFullL2),
        .PCL_wbHold(                        PCL_wbHold),
        .PCL_wbStorageEnd(                  PCL_wbStorageEnd),
        .PCL_wbStorageOp(                   PCL_wbStorageOp),
        .PGM_apuPresent(                    PGM_coprocPresent),
        .TRC_fifoFull(                      TRC_fifoFull),
        .TRC_fifoOneEntryFree(              TRC_fifoOneEntryFree),
        .TRC_se(                            TRC_se),
        .TRC_seCtrEqZeroL2(                 TRC_seCtrEqZeroL2),
        .TRC_sleepReq(                      TRC_sleepReq),
        .VCT_anySwap(                       VCT_anySwap),
        .VCT_msrWE(                         VCT_msrWEL2),
        .VCT_swap01(                        VCT_swap01),
        .VCT_swap23(                        VCT_swap23),
        .VCT_vectorBus(                     VCT_vectorBus[0:7]),
        .VCT_wbFlush(                       VCT_wbFlush),
        .VCT_wbRfci(                        VCT_wbRfci),
        .VCT_wbRfi(                         VCT_wbRfi),
        .VCT_wbSuppress(                    VCT_wbSuppress),
        .XXX_traceDisable(                  TRC_c405TraceDisable),
        .coreReset(                         resetCore),
        .dcdValidOp_Neg(                    dcdApuValidOp_NEG),
        .MMU_isParityErr(                   MMU_isParityErr),
        .ICU_parityErrE(                    ICU_parityErrE),
        .ICU_parityErrO(                    ICU_parityErrO),
        .ICU_tagParityErr(                  ICU_tagParityErr),
        .IFB_exeISideMachChk(               IFB_exeISideMachChk),
        .ICU_CCR0IPE(                       ICU_CCR0IPE),
        .ICU_CCR0TPE(                       ICU_CCR0TPE)
        );

p405s_exe_top
 exe_topSch(
        .EXE_admMco(                        EXE_admMco),
        .EXE_apuLoadData(                   EXE_apuLoadData[0:31]),
        .EXE_cc(                            EXE_cc[0:3]),
        .EXE_dac1CO(                        EXE_dac1GtDsEa),
        .EXE_dac1SumBit30Eq(                EXE_dac1Bits30Eq),
        .EXE_dac1SumBit31Eq(                EXE_dac1Bits31Eq),
        .EXE_dac1SumBits0thru27Eq(          EXE_dac1Bits0to26Eq),
        .EXE_dac1SumBits28and29Eq(          EXE_dac1Bits27to29Eq),
        .EXE_dac2CO(                        EXE_dac2GtDsEa),
        .EXE_dac2SumBit30Eq(                EXE_dac2Bits30Eq),
        .EXE_dac2SumBit31Eq(                EXE_dac2Bits31Eq),
        .EXE_dac2SumBits0thru27Eq(          EXE_dac2Bits0to26Eq),
        .EXE_dac2SumBits28and29Eq(          EXE_dac2Bits27to29Eq),
        .EXE_dcrAddr(                       EXE_dcrAddr[0:9]),
        .EXE_dcrDataBus(                    EXE_dcrDataBus[0:31]),
        .EXE_dcuData(                       EXE_dcuData[0:31]),
        .EXE_divMco(                        EXE_divMco),
        .EXE_dofDregParityErrL2(            EXE_dofDregParityErrL2),
        .EXE_dsEA_NEG(                      EXE_dsEA_NEG[0:31]),
        .EXE_dsEaCP_NEG(                    EXE_dsEaCP[0:7]),
        .EXE_dvc1ByteCmp(                   EXE_dvc1ByteCmp[0:3]),
        .EXE_dvc2ByteCmp(                   EXE_dvc2ByteCmp[0:3]),
        .EXE_ea(                            EXE_ea[30:31]),
        .EXE_eaARegBuf(                     EXE_eaARegBuf[0:21]),
        .EXE_eaBRegBuf(                     EXE_eaBRegBuf[0:21]),
        .EXE_ifbSprDataBus(                 EXE_ifbSprDataBus[0:31]),
        .EXE_mmuIcuSprDataBus(              EXE_mmuIcuSprDataBus[0:31]),
        .EXE_multMco(                       EXE_multMco),
        .EXE_raData(                        EXE_raData[0:31]),
        .EXE_rbData(                        EXE_rbData[0:31]),
        .EXE_sprAddr(                       EXE_sprAddr[4:9]),
        .EXE_timJtgSprDataBus(              EXE_timJtgSprDataBus[0:31]),
        .EXE_trap(                          EXE_trap),
        .EXE_vctDbgSprDataBus(              EXE_vctDbgSprDataBus[0:31]),
        .EXE_wrteeIn(                       EXE_wrteeIn),
        .EXE_xer(                           EXE_xer[0:2]),
        .EXE_xerCa(                         EXE_xerCa),
        .EXE_xerTBC(                        EXE_xerTBC[0:6]),
        .EXE_xerTBCIn(                      EXE_xerTBCIn[0:6]),
        .EXE_xerTBCNotEqZero(               EXE_xerTBCNotEqZero),
        .APU_exeCa(                         APU_exeCa),
        .APU_exeCr(                         APU_exeCr[0:3]),
        .APU_exeOv(                         APU_exeOv),
        .APU_exeResult(                     APU_exeResult[0:31]),
        .CB(                                CB),
        .DBG_dacEn(                         DBG_dacEn),
        .DBG_sprDataBus(                    DBG_sprDataBus[0:31]),
        .DCU_SDQ_mod_NEG(                   DCU_SDQ_mod[0:31]),
        .DCU_data_NEG(                      DCU_data_NEG[0:31]),
        .DCU_parityError(                   DCU_parityError),
        .ICU_sprDataBus(                    ICU_sprDataBus[0:31]),
        .IFB_exeMcrxr(                      IFB_exeMcrxrL2),
        .IFB_exeOpForExe2L2(                IFB_exeOpForExe2L2),
        .IFB_sprDataBus(                    IFB_sprDataBus[0:31]),
        .JTG_sprDataBus(                    JTG_sprDataBus[0:31]),
        .LSSD_coreTestEn(                   LSSD_coreTestEn),
        .MMU_sprDataBus(                    MMU_sprDataBus[0:31]),
        .OCM_dsData(                        OCM_dsData[0:31]),
        .PCL_aPortRregBypass(               PCL_aPortRregBypass),
        .PCL_aRegE2(                        PCL_aRegG2),
        .PCL_aRegForEaE2(                   PCL_aRegForEaE2),
        .PCL_abRegE1(                       PCL_aRegG1),
        .PCL_addFour(                       PCL_addFour),
        .PCL_apuTrcLoadEn(                  PCL_apuLoadEn),
        .PCL_bPortLitGenSel(                PCL_bPortLitGenSel),
        .PCL_bPortRregBypass(               PCL_bPortRregBypass),
        .PCL_bRegE2(                        PCL_bRegG2),
        .PCL_bRegForEaE2(                   PCL_bRegForEaE2),
        .PCL_dRegBypassMuxSel(              PCL_dRegBypassMuxSel),
        .PCL_dRegE1(                        PCL_dRegE1),
        .PCL_dbgSprDcds(                    PCL_dbgSprDcds[0:3]),
        .PCL_dcdApAddr(                     PCL_dcdApAddr[0:9]),
        .PCL_dcdAregLoadUse(                PCL_aPortDcdLoadUse),
        .PCL_dcdBpAddr(                     PCL_dcdBpAddr[0:9]),
        .PCL_dcdBregLoadUse(                PCL_bPortDcdLoadUse),
        .PCL_dcdHotCIn(                     PCL_dcdHotCIn),
        .PCL_dcdImmd(                       PCL_dcdImmd[11:31]),
        .PCL_dcdLitCntl(                    PCL_dcdLitCntl[0:4]),
        .PCL_dcdMdSelQ(                     PCL_dcdMdSel),
        .PCL_dcdMrSelQ(                     PCL_dcdMrSel),
        .PCL_dcdSpAddr(                     PCL_dcdSpAddr[0:9]),
        .PCL_dcdSregLoadUse(                PCL_sPortDcdLoadUse),
        .PCL_dcdSrmBpSel(                   PCL_dcdSrmMuxSel[0:2]),
        .PCL_dcdXerCa(                      PCL_dcdXerCa),
        .PCL_dofDregE1(                     PCL_dofDregE1),
        .PCL_dofDregMuxSel(                 PCL_dofDregMuxSel[0:1]),
        .PCL_dvcByteEnL2(                   PCL_dvcByteEnL2[0:3]),
        .PCL_dvcCmpEn(                      PCL_dvcCmpEn),
        .PCL_exe2AccRegMuxSel(              PCL_exe2AccRegMuxSel[0:1]),
        .PCL_exe2Hold(                      PCL_exe2Hold),
        .PCL_exe2MacEn(                     PCL_exe2MacEn),
        .PCL_exe2MacOrMultEnForMS(          PCL_exe2MacOrMultEnForMS[0:1]),
        .PCL_exe2MacOrMultEn_NEG(           PCL_exe2MacOrMultEn_NEG[0:1]),
        .PCL_exe2MacSat(                    PCL_exe2MacSat),
        .PCL_exe2MultEn(                    PCL_exe2MultEn),
        .PCL_exe2MultHiWd(                  PCL_exe2MultHiWd),
        .PCL_exe2NegMac(                    PCL_exe2NegMac),
        .PCL_exe2SignedOp(                  PCL_exe2SignedOp),
        .PCL_exe2XerOvEn(                   PCL_exe2XerOvEn),
        .PCL_exeAddEn(                      PCL_exeAddEn),
        .PCL_exeAddSgndOp_NEG(              PCL_exeAddSgndOp_NEG[0:1]),
        .PCL_exeAdmCntl(                    PCL_exeAdmCntl[0:3]),
        .PCL_exeApuValidOp(                 PCL_exeValidOp),
        .PCL_exeAregLoadUse(                PCL_aPortExeLoadUse),
        .PCL_exeBregLoadUse(                PCL_bPortExeLoadUse),
        .PCL_exeCmplmntA(                   PCL_exeCmplmntA),
        .PCL_exeCmplmntA_NEG(               PCL_exeCmplmntA_NEG),
        .PCL_exeDivEn(                      PCL_exeDivEn),
        .PCL_exeDivEnForLSSD(               PCL_exeDivEnForLSSD),
        .PCL_exeDivEnForMuxSel(             PCL_exeDivEnForMuxSel[0:1]),
        .PCL_exeDivEn_NEG(                  PCL_exeDivEn_NEG),
        .PCL_exeDivSgndOp(                  PCL_exeDivSgndOp),
        .PCL_exeDvcHold(                    PCL_exeDvcHold),
        .PCL_exeEaCalc(                     PCL_exeEaCalc),
        .PCL_exeEaQwEn(                     PCL_exeEaQwEn[0:3]),
        .PCL_exeFpuOp(                      PCL_exeFpuOp),
        .PCL_exeLoadUseHold(                PCL_exeLoadUseHold),
        .PCL_exeLogicalCntl(                PCL_exeLogicalCntl[0:7]),
        .PCL_exeLogicalUnitEnForLSSD(       PCL_exeLogicalUnitEnForLSSD),
        .PCL_exeLogicalUnitEn_NEG(          PCL_exeLogicalUnitEn),
        .PCL_exeMacEn(                      PCL_exeMacEn),
        .PCL_exeMacOrMultEn_NEG(            PCL_exeMacOrMultEn),
        .PCL_exeMfspr(                      PCL_mfSPR),
        .PCL_exeMtspr(                      PCL_mtSPR),
        .PCL_exeMultEn(                     PCL_exeMultEn),
        .PCL_exeMultEnForMuxSel(            PCL_exeMultEnForMuxSel[0:1]),
        .PCL_exeMultEn_NEG(                 PCL_exeMultEn_NEG[0:1]),
        .PCL_exeNegMac(                     PCL_exeexeNegMac),
        .PCL_exeRaEn(                       PCL_exeRaEn[0:3]),
        .PCL_exeRbEn(                       PCL_exeRbEn[0:3]),
        .PCL_exeSprDataEn_NEG(              PCL_exeSprDataEn),
        .PCL_exeSprDcds(                    PCL_exeSprDcds[0:4]),
        .PCL_exeSprUnitEn_NEG(              PCL_exeSprUnitEn),
        .PCL_exeSregLoadUse(                PCL_sPortExeLoadUse),
        .PCL_exeSrmBpSel(                   PCL_exeSrmBpSel[0:2]),
        .PCL_exeSrmCntl(                    PCL_exeSrmCntl[0:3]),
        .PCL_exeSrmUnitEnForLSSD(           PCL_exeSrmUnitEnForLSSD),
        .PCL_exeSrmUnitEn_NEG(              PCL_exeSrmUnitEn),
        .PCL_exeTrapCond(                   PCL_exeTrapCond[0:4]),
        .PCL_exeWrtee(                      PCL_exeWrtee),
        .PCL_exeXerCaEn(                    PCL_exeXerCaEn),
        .PCL_exeXerOvEn(                    PCL_exeXerOvEn),
        .PCL_gateZeroToAreg(                PCL_gateZeroToAreg),
        .PCL_gateZeroToSreg(                PCL_gateZeroToSreg),
        .PCL_holdCIn(                       PCL_holdCIn),
        .PCL_holdMdMr(                      PCL_holdMdMr),
        .PCL_ldAdjE1(                       PCL_ldAdjE1),
        .PCL_ldAdjE2(                       PCL_ldAdjG1[1:3]),
        .PCL_ldAdjMuxSel(                   PCL_ldAdjMuxSel[0:1]),
        .PCL_ldFillByPassMuxSel(            PCL_ldFillByPassMuxSel[0:5]),
        .PCL_ldMuxSel(                      PCL_ldMuxSel[0:7]),
        .PCL_ldSteerMuxSel(                 PCL_ldSteerMuxSel[0:7]),
        .PCL_lwbLpAddr(                     PCL_lwbLpAddr[0:4]),
        .PCL_lwbLpEqdcdApAddr(              PCL_LpEqAp),
        .PCL_lwbLpEqdcdBpAddr(              PCL_LpEqBp),
        .PCL_lwbLpEqdcdSpAddr(              PCL_LpEqSp),
        .PCL_lwbLpWrEn(                     PCL_lwbLpWE),
        .PCL_mfDCRL2(                       PCL_mfDCRL2),
        .PCL_resultMuxSel(                  PCL_resultMuxSel),
        .PCL_resultRegE1(                   PCL_resultRegG1),
        .PCL_resultRegE2(                   PCL_resultRegG2),
        .PCL_sPortRregBypass(               PCL_sPortRregBypass),
        .PCL_sRegE1(                        PCL_sRegG1),
        .PCL_sRegE2(                        PCL_sRegG2),
        .PCL_sdqMuxSel(                     PCL_sdqMuxSel),
        .PCL_sprHold(                       PCL_ifbSprHold),
        .PCL_sraRegE1(                      PCL_sraRegG1),
        .PCL_sraRegE2(                      PCL_sraRegE2),
        .PCL_srmRegE1(                      PCL_srmRegG1),
        .PCL_srmRegE2(                      PCL_srmRegE2[0:2]),
        .PCL_timSprDcds(                    PCL_timSprDcds[0:5]),
        .PCL_vctSprDcds(                    PCL_vctSprDcds[0:5]),
        .PCL_wbHold(                        PCL_wbHold),
        .PCL_wbRpAddr(                      PCL_wbRpAddr[0:4]),
        .PCL_wbRpEqdcdApAddr(               PCL_RpEqAp),
        .PCL_wbRpEqdcdBpAddr(               PCL_RpEqBp),
        .PCL_wbRpEqdcdSpAddr(               PCL_RpEqSp),
        .PCL_wbRpWrEn(                      PCL_wbRpWE),
        .PCL_xerL2Hold(                     PCL_xerL2Hold),
        .PGM_deterministicMult(             PGM_deterministicMult),
        .TIM_sprDataBus(                    TIM_sprDataBus[0:31]),
        .VCT_sprDataBus(                    VCT_sprDataBus[0:31]),
        .XXX_dcrDataBus(                    XXX_dcrDataBus[0:31]),
        .PCL_exeDvcOrParityHold(            PCL_exeDvcOrParityHold),
        .coreReset(                         resetCore),
        .PCL_BpEqSp(                        PCL_BpEqSp),
	      .EXE_gprSysClkPI(                   EXE_gprSysClkPI),
 	      .EXE_gprRen(                        PCL_gprRdClk)
        );

p405s_pcl_top
 pcl_topSch(
        .PCL_LpEqSp(                        PCL_LpEqSp),
        .PCL_Rbit(                          PCL_Rbit),
        .PCL_aPortRregBypass(               PCL_aPortRregBypass),
        .PCL_aRegE2(                        PCL_aRegG2),
        .PCL_aRegForEaE2(                   PCL_aRegForEaE2),
        .PCL_abRegE1(                       PCL_aRegG1),
        .PCL_addFour(                       PCL_addFour),
        .PCL_apuDcdHold(                    PCL_dcdHoldForApu),
        .PCL_apuExeFlush(                   PCL_exeFlushForApu),
        .PCL_apuExeHold(                    PCL_exeHoldForApu),
        .PCL_apuExeWdCnt(                   PCL_apuExeWdCnt[0:1]),
        .PCL_apuLwbLoadDV(                  PCL_apuLoadDV),
        .PCL_apuTrcLoadEn(                  PCL_apuLoadEn),
        .PCL_apuWbHold(                     PCL_apuWbHold),
        .PCL_bPortLitGenSel(                PCL_bPortLitGenSel),
        .PCL_bPortRregBypass(               PCL_bPortRregBypass),
        .PCL_bRegE2(                        PCL_bRegG2),
        .PCL_bRegForEaE2(                   PCL_bRegForEaE2),
        .PCL_blkFlush(                      PCL_blkFlush),
        .PCL_blkFlushForVct(                PCL_blkFlushForVct[0:2]),
        .PCL_dIcmpForStep(                  PCL_dIcmpForStep),
        .PCL_dIcmpForStuff(                 PCL_dIcmpForStuff),
        .PCL_dIcmpForWbFlushQDlydL2(        PCL_dIcmpForWbFlushQDlydL2),
        .PCL_dRegBypassMuxSel(              PCL_dRegBypassMuxSel),
        .PCL_dRegE1(                        PCL_dRegE1),
        .PCL_dbgSprDcds(                    PCL_dbgSprDcds[0:3]),
        .PCL_dcdApAddr(                     PCL_dcdApAddr[0:9]),
        .PCL_dcdAregLoadUse(                PCL_aPortDcdLoadUse),
        .PCL_dcdBpAddr(                     PCL_dcdBpAddr[0:9]),
        .PCL_dcdBregLoadUse(                PCL_bPortDcdLoadUse),
        .PCL_dcdHoldForIfb(                 PCL_dcdHoldForIfb[0:2]),
        .PCL_dcdHotCIn(                     PCL_dcdHotCIn),
        .PCL_dcdImmd(                       PCL_dcdImmd[11:31]),
        .PCL_dcdLitCntl(                    PCL_dcdLitCntl[0:4]),
        .PCL_dcdMdSelQ(                     PCL_dcdMdSel),
        .PCL_dcdMrSelQ(                     PCL_dcdMrSel),
        .PCL_dcdSpAddr(                     PCL_dcdSpAddr[0:9]),
        .PCL_dcdSregLoadUse(                PCL_sPortDcdLoadUse),
        .PCL_dcdSrmBpSel(                   PCL_dcdSrmMuxSel[0:2]),
        .PCL_dcdXerCa(                      PCL_dcdXerCa),
        .PCL_dcuByteEn(                     PCL_dcuByteEn[0:3]),
        .PCL_dcuOp(                         PCL_dcuOp[0:11]),
        .PCL_dcuOp_early(                   PCL_dcuOp_early[0:2]),
        .PCL_diagBus(                       PCL_diagBus[0:9]),
        .PCL_dofDRegE1(                     PCL_dofDregE1),
        .PCL_dofDregFull(                   PCL_dofDregFull),
        .PCL_dofDRegMuxSel(                 PCL_dofDregMuxSel[0:1]),
        .PCL_dsMmuOp(                       PCL_dsMmuOp[0:3]),
        .PCL_dsOcmByteEn(                   PCL_dsOcmByteEn[0:3]),
        .PCL_dvcByteEnL2(                   PCL_dvcByteEnL2[0:3]),
        .PCL_dvcCmpEn(                      PCL_dvcCmpEn),
        .PCL_exe2AccRegMuxSel(              PCL_exe2AccRegMuxSel[0:1]),
        .PCL_exe2ClearOrFlush(              PCL_exe2FlushorClear),
        .PCL_exe2DataE1(                    PCL_exe2DataE1),
        .PCL_exe2DataE2(                    PCL_exe2DataE2),
        .PCL_exe2Full(                      PCL_exe2Full),
        .PCL_exe2Hold(                      PCL_exe2Hold),
        .PCL_exe2IarE1(                     PCL_exe2IarE1),
        .PCL_exe2IarE2(                     PCL_exe2IarE2),
        .PCL_exe2MacEn(                     PCL_exe2MacEn),
        .PCL_exe2MacOrMultEnForMS(          PCL_exe2MacOrMultEnForMS[0:1]),
        .PCL_exe2MacOrMultEn_NEG(           PCL_exe2MacOrMultEn_NEG[0:1]),
        .PCL_exe2MacSat(                    PCL_exe2MacSat),
        .PCL_exe2MultEn(                    PCL_exe2MultEn),
        .PCL_exe2MultHiWd(                  PCL_exe2MultHiWd),
        .PCL_exe2NegMac(                    PCL_exe2NegMac),
        .PCL_exe2SignedOp(                  PCL_exe2SignedOp),
        .PCL_exe2XerOvEn(                   PCL_exe2XerOvEn),
        .PCL_exeAbort(                      PCL_exeAbort),
        .PCL_exeAddEn(                      PCL_exeAddEn),
        .PCL_exeAddSgndOp_NEG(              PCL_exeAddSgndOp_NEG[0:1]),
        .PCL_exeAdmCntl(                    PCL_exeAdmCntl[0:3]),
        .PCL_exeApuOp(                      PCL_exeApuOp),
        .PCL_exeApuValidOp(                 PCL_exeValidOp),
        .PCL_exeAregLoadUse(                PCL_aPortExeLoadUse),
        .PCL_exeBregLoadUse(                PCL_bPortExeLoadUse),
        .PCL_exeCmplmntA(                   PCL_exeCmplmntA),
        .PCL_exeCmplmntA_NEG(               PCL_exeCmplmntA_NEG),
        .PCL_exeCpuOp(                      PCL_exeIllegalOpLtch),
        .PCL_exeDbgLdOp(                    PCL_exeDbgLdOp),
        .PCL_exeDbgRdOp(                    PCL_exeDbgRdOp),
        .PCL_exeDbgStOp(                    PCL_exeDbgStOp),
        .PCL_exeDbgWrOp(                    PCL_exeDbgWrOp),
        .PCL_exeDivEn(                      PCL_exeDivEn),
        .PCL_exeDivEnForLSSD(               PCL_exeDivEnForLSSD),
        .PCL_exeDivEnForMuxSel(             PCL_exeDivEnForMuxSel[0:1]),
        .PCL_exeDivEn_NEG(                  PCL_exeDivEn_NEG),
        .PCL_exeDivSgndOp(                  PCL_exeDivSgndOp),
        .PCL_exeDvcHold(                    PCL_exeDvcHold),
        .PCL_exeDvcOrParityHold(            PCL_exeDvcOrParityHold),
        .PCL_exeEaCalc(                     PCL_exeEaCalc),
        .PCL_exeEaQwEn(                     PCL_exeEaQwEn[0:3]),
        .PCL_exeFpuOp(                      PCL_exeFpuOp),
        .PCL_exeFull(                       PCL_exeFull),
        .PCL_exeHoldForCr(                  PCL_exeHoldForCr),
        .PCL_exeIarHold(                    PCL_exeIarHold),
        .PCL_exeLdNotSt(                    PCL_exeLdNotSt),
        .PCL_exeLoadUseHold(                PCL_exeLoadUseHold),
        .PCL_exeLogicalCntl(                PCL_exeLogicalCntl[0:7]),
        .PCL_exeLogicalUnitEnForLSSD(       PCL_exeLogicalUnitEnForLSSD),
        .PCL_exeLogicalUnitEn_NEG(          PCL_exeLogicalUnitEn),
        .PCL_exeMacEn(                      PCL_exeMacEn),
        .PCL_exeMacOrMultEn_NEG(            PCL_exeMacOrMultEn),
        .PCL_exeMultEn(                     PCL_exeMultEn),
        .PCL_exeMultEnForMuxSel(            PCL_exeMultEnForMuxSel[0:1]),
        .PCL_exeMultEn_NEG(                 PCL_exeMultEn_NEG[0:1]),
        .PCL_exeNegMac(                     PCL_exeexeNegMac),
        .PCL_exePrivOp(                     PCL_exePrivOp),
        .PCL_exeRaEn(                       PCL_exeRaEn[0:3]),
        .PCL_exeRbEn(                       PCL_exeRbEn[0:3]),
        .PCL_exeSprDataEn_NEG(              PCL_exeSprDataEn),
        .PCL_exeSprDcds(                    PCL_exeSprDcds[0:4]),
        .PCL_exeSprUnitEn_NEG(              PCL_exeSprUnitEn),
        .PCL_exeSregLoadUse(                PCL_sPortExeLoadUse),
        .PCL_exeSrmBpSel(                   PCL_exeSrmBpSel[0:2]),
        .PCL_exeSrmCntl(                    PCL_exeSrmCntl[0:3]),
        .PCL_exeSrmUnitEnForLSSD(           PCL_exeSrmUnitEnForLSSD),
        .PCL_exeSrmUnitEn_NEG(              PCL_exeSrmUnitEn),
        .PCL_exeStorageOp(                  PCL_exeStorageOp),
        .PCL_exeStringMultiple(             PCL_exeStringMultiple),
        .PCL_exeTlbOp(                      PCL_exeTlbOp),
        .PCL_exeTrap(                       PCL_exeTrap),
        .PCL_exeTrapCond(                   PCL_exeTrapCond[0:4]),
        .PCL_exeWrExtEn(                    PCL_exeWrExtEn),
        .PCL_exeWrtee(                      PCL_exeWrtee),
        .PCL_exeXerCaEn(                    PCL_exeXerCaEn),
        .PCL_exeXerOvEn(                    PCL_exeXerOvEn),
        .PCL_gateZeroToAreg(                PCL_gateZeroToAreg),
        .PCL_gateZeroToSreg(                PCL_gateZeroToSreg),
        .PCL_holdCIn(                       PCL_holdCIn),
        .PCL_holdMdMr(                      PCL_holdMdMr),
        .PCL_icuOp(                         PCL_icuOp[0:3]),
        .PCL_icuSprDcds(                    EXE_icuSprDcds[0:2]),
        .PCL_ifbSprHold(                    PCL_ifbSprHold),
        .PCL_jtgSprDcd(                     PCL_jtgSprDcd),
        .PCL_ldAdjE1(                       PCL_ldAdjE1),
        .PCL_ldAdjE2(                       PCL_ldAdjG1[1:3]),
        .PCL_ldAdjMuxSel(                   PCL_ldAdjMuxSel[0:1]),
        .PCL_ldFillBypassMuxSel(            PCL_ldFillByPassMuxSel[0:5]),
        .PCL_ldMuxSel(                      PCL_ldMuxSel[0:7]),
        .PCL_ldSteerMuxSel(                 PCL_ldSteerMuxSel[0:7]),
        .PCL_lwbCacheableL2(                PCL_lwbCacheableL2),
        .PCL_lwbLpAddr(                     PCL_lwbLpAddr[0:4]),
        .PCL_lwbLpEqdcdApAddr(              PCL_LpEqAp),
        .PCL_lwbLpEqdcdBpAddr(              PCL_LpEqBp),
        .PCL_lwbLpWrEn(                     PCL_lwbLpWE),
        .PCL_mfDCR(                         PCL_mfDCR),
        .PCL_mfDCRL2(                       PCL_mfDCRL2),
        .PCL_mfSPR(                         PCL_mfSPR),
        .PCL_mmuExeAbort(                   PCL_mmuExeAbort),
        .PCL_mmuIcuSprHold(                 PCL_mmuIcuSprHold),
        .PCL_mmuSprDcd(                     PCL_mmuSprDcd[0:8]),
        .PCL_mtDCR(                         PCL_mtDCR),
        .PCL_mtSPR(                         PCL_mtSPR),
        .PCL_ocmAbortReq(                   PCL_ocmAbortReq),
        .PCL_resultMuxSel(                  PCL_resultMuxSel),
        .PCL_resultRegE1(                   PCL_resultRegG1),
        .PCL_resultRegE2(                   PCL_resultRegG2),
        .PCL_sPortRregBypass(               PCL_sPortRregBypass),
        .PCL_sRegE1(                        PCL_sRegG1),
        .PCL_sRegE2(                        PCL_sRegG2),
        .PCL_sdqMuxSel(                     PCL_sdqMuxSel),
        .PCL_sraRegE1(                      PCL_sraRegG1),
        .PCL_sraRegE2(                      PCL_sraRegE2),
        .PCL_srmRegE1(                      PCL_srmRegG1),
        .PCL_srmRegE2(                      PCL_srmRegE2[0:2]),
        .PCL_stSteerCntl(                   PCL_stSteerCntl[0:9]),
        .PCL_timJtgSprHold(                 PCL_timJtgsprHold),
        .PCL_timSprDcds(                    PCL_timSprDcds[0:5]),
        .PCL_tlbRE(                         PCL_tlbRE),
        .PCL_tlbSX(                         PCL_tlbSX),
        .PCL_tlbWE(                         PCL_tlbWE),
        .PCL_tlbWS(                         PCL_tlbWS),
        .PCL_trcLoadDV(                     PCL_trcLoadDV),
        .PCL_vctDbgSprHold(                 PCL_vctDbgsprHold),
        .PCL_vctSprDcds(                    PCL_vctSprDcds[0:5]),
        .PCL_wbAlgnErr(                     PCL_algnErr),
        .PCL_wbClearOrFlush(                PCL_wbClear),
        .PCL_wbClearTerms(                  PCL_wbClearTerms),
        .PCL_wbComplete(                    PCL_wbComplete),
        .PCL_wbDbgIcmp(                     PCL_wbDbgIcmp),
        .PCL_wbFullForPO(                   PCL_wbFull),
        .PCL_wbFullL2(                      PCL_wbFullL2),
        .PCL_wbHold(                        PCL_wbHold),
        .PCL_wbHoldNonErr(                  PCL_wbHoldNonErr),
        .PCL_wbLdNotSt(                     PCL_wbLdNotSt),
        .PCL_wbRpAddr(                      PCL_wbRpAddr[0:4]),
        .PCL_wbRpEqdcdApAddr(               PCL_RpEqAp),
        .PCL_wbRpEqdcdBpAddr(               PCL_RpEqBp),
        .PCL_wbRpEqdcdSpAddr(               PCL_RpEqSp),
        .PCL_wbRpWrEn(                      PCL_wbRpWE),
        .PCL_wbStorageOp(                   PCL_wbStorageOp),
        .PCL_wbStrgEnd(                     PCL_wbStorageEnd),
        .PCL_xerL2Hold(                     PCL_xerL2Hold),
        .APU_dcdApuOp(                      APU_dcdApuOp),
        .APU_dcdExeLdDepend(                APU_dcdExeLdDepend),
        .APU_dcdForceAlgn(                  APU_dcdForceAlgn),
        .APU_dcdForceBESteering(            APU_dcdForceBESteering),
        .APU_dcdFpuOp(                      APU_dcdFpuOp),
        .APU_dcdGprWr(                      APU_dcdGprWr),
        .APU_dcdLdStByte(                   APU_dcdLdStByte),
        .APU_dcdLdStDw(                     APU_dcdLdStDw),
        .APU_dcdLdStHw(                     APU_dcdLdStHw),
        .APU_dcdLdStQw(                     APU_dcdLdStQw),
        .APU_dcdLdStWd(                     APU_dcdLdStWd),
        .APU_dcdLoad(                       APU_dcdLoad),
        .APU_dcdLwbLdDepend(                APU_dcdLwbLdDepend),
        .APU_dcdPrivOp(                     APU_dcdPrivOp),
        .APU_dcdRaEn(                       APU_dcdRaEn),
        .APU_dcdRbEn(                       APU_dcdRbEn),
        .APU_dcdStore(                      APU_dcdStore),
        .APU_dcdTrapBE(                     APU_dcdTrapBE),
        .APU_dcdTrapLE(                     APU_dcdTrapLE),
        .APU_dcdUpdate(                     APU_dcdUpdate),
        .APU_dcdWbLdDepend(                 APU_dcdWbLdDepend),
        .APU_dcdXerCAEn(                    APU_dcdXerCAEn),
        .APU_dcdXerOVEn(                    APU_dcdXerOVEn),
        .APU_exeBlkingMco(                  APU_exeBlkingMco),
        .APU_exeBusy(                       APU_exeBusy),
        .APU_exeNonBlkingMco(               APU_exeNonBlkingMco),
        .CAR_cacheable(                     CAR_cacheable),
        .CAR_endian(                        CAR_endian),
        .CB(                                CB),
        .DBG_dvcRdEn(                       DBG_dvcRdEn),
        .DBG_dvcWrEn(                       DBG_dvcWrEn),
        .DBG_exeIacSuppress(                DBG_exeIacSuppress),
        .DBG_icmpEn(                        DBG_icmpEn),
        .DBG_wbDacSuppress(                 DBG_wbDacSuppress),
        .DCU_CA(                            DCU_CA),
        .DCU_DA(                            DCU_DA),
        .DCU_DOF(                           PGM_dcu_DOF),
        .DCU_carByteEn(                     DCU_carByteEn[0:3]),
        .DCU_firstCycCarStXltV(             DCU_firstCycCarStXltV),
        .DCU_pclOcmLdPendNoWait(            DCU_pclOcmWait),
        .EXE_admMco(                        EXE_admMco),
        .EXE_divMco(                        EXE_divMco),
        .EXE_ea(                            EXE_ea[30:31]),
        .EXE_multMco(                       EXE_multMco),
        .EXE_trap(                          EXE_trap),
        .EXE_xerTBC(                        EXE_xerTBC[0:6]),
        .EXE_xerTBCIn(                      EXE_xerTBCIn[0:6]),
        .EXE_xerTBCNotEqZero(               EXE_xerTBCNotEqZero),
        .ICU_CCR0DPP(                       ICU_CCR0DPP),
        .ICU_LDBE(                          ICU_LDBE),
        .ICU_dsCA(                          ICU_dsCA),
        .ICU_gprDRCC(                       ICU_GPRC),
        .IFB_dcdBubble(                     IFB_dcdBubble),
        .IFB_dcdDataIn_NEG(                 IFB_dcdDataIn_Neg[0:31]),
        .IFB_dcdFull(                       IFB_dcdFullL2[0]),
        .IFB_dcdRegE1(                      IFB_dcdRegE1),
        .IFB_dcdRegE2(                      IFB_dcdRegE2),
        .IFB_exeCorrect(                    IFB_exeCorrect),
        .IFB_exeFlush(                      IFB_exeFlushB),
        .IFB_exeRfciL2(                     IFB_exeRfciL2),
        .IFB_exeRfiL2(                      IFB_exeRfiL2),
        .IFB_exeScL2(                       IFB_exeScL2),
        .IFB_stepStL2(                      IFB_stepStL2),
        .IFB_stuffStL2(                     IFB_stuffStL2),
        .IFB_trcPipeHold(                   IFB_tracePipeHold),
        .LSSD_coreTestEn(                   LSSD_coreTestEn),
        .MMU_BMCO(                          MMU_BMCO),
        .MMU_dsStatus(                      MMU_dsStatus[0:4]),
        .MMU_wbHold(                        MMU_wbHold),
        .OCM_DOF(                           OCM_DOF),
        .OCM_dsComplete(                    OCM_dsComplete),
        .PGM_divEn(                         PGM_divEn),
        .PGM_mmuEn(                         PGM_mmuEn),
        .VCT_errorSprSuppress(              VCT_errorSprSuppress),
        .VCT_exeSuppForApu(                 VCT_exeSuppForApu),
        .VCT_exeSuppForCr(                  VCT_exeSuppForCr),
        .VCT_exeSuppForExe2Clear(           VCT_exeSuppForExe2Clear),
        .VCT_exeSuppress(                   VCT_exeSuppress),
        .VCT_sxrOR_L2(                      VCTsxrOR_L2),
        .VCT_wbFlush(                       VCT_wbFlush),
        .VCT_wbFlushAsync(                  VCT_wbFlushAsync),
        .VCT_wbLoadSuppress(                VCT_wbLoadSuppress),
        .VCT_wbSuppress(                    VCT_wbSuppress),
        .XXX_dcrAck(                        XXX_dcrAck),
        .c2Clk(                             c2Clk),
        .coreReset(                         resetCore),
        .dcdApuValidOp_NEG(                 dcdApuValidOp_NEG),
        .lwbFullL2(                         lwbFullL2),
        .PCL_BpEqSp                        (PCL_BpEqSp),
	.PCL_gprRdClk                      (PCL_gprRdClk)
        );

endmodule
