library verilog;
use verilog.vl_types.all;
entity p405s_fetcherCntl is
    port(
        IFB_TEL2        : out    vl_logic;
        IFB_TETypeL2    : out    vl_logic_vector(0 to 10);
        IFB_cntxSync    : out    vl_logic;
        IFB_cntxSyncOCM : out    vl_logic;
        IFB_coreSleepReqL2: out    vl_logic;
        IFB_dcdFullApuL2: out    vl_logic;
        IFB_dcdFullL2   : out    vl_logic_vector(0 to 1);
        IFB_diagBus     : out    vl_logic_vector(0 to 7);
        IFB_exeFlushA   : out    vl_logic;
        IFB_exeFlushB   : out    vl_logic;
        IFB_extStopAck  : out    vl_logic;
        IFB_fetchReq    : out    vl_logic;
        IFB_icuCancelDataL2: out    vl_logic;
        IFB_isAbortForICU: out    vl_logic_vector(0 to 2);
        IFB_isAbortForMMU: out    vl_logic;
        IFB_nonSpecAcc  : out    vl_logic;
        IFB_ocmAbort    : out    vl_logic;
        IFB_postEntry   : out    vl_logic;
        IFB_rstStepPend : out    vl_logic;
        IFB_rstStuffPend: out    vl_logic;
        IFB_stopAck     : out    vl_logic;
        IFB_traceESL2   : out    vl_logic_vector(0 to 1);
        IFB_traceType   : out    vl_logic_vector(0 to 1);
        coreResetL2     : out    vl_logic;
        dbdrPulseCntlE1 : out    vl_logic;
        dcdApuE1        : out    vl_logic;
        dcdBrTarSel     : out    vl_logic_vector(0 to 1);
        dcdBubble       : out    vl_logic;
        dcdClear        : out    vl_logic;
        dcdDataMuxSel   : out    vl_logic_vector(0 to 1);
        dcdE1           : out    vl_logic;
        dcdE2           : out    vl_logic;
        dcdFlush        : out    vl_logic;
        dcdFullL2       : out    vl_logic;
        dcdIarMuxSel    : out    vl_logic_vector(0 to 1);
        exeClear        : out    vl_logic;
        exeDataE1       : out    vl_logic;
        exeDataE2       : out    vl_logic;
        exeDataSel      : out    vl_logic;
        exeFlush        : out    vl_logic;
        exeFlushorClear : out    vl_logic;
        exeFullL2       : out    vl_logic;
        exeIarE2        : out    vl_logic;
        isEA_22DlyL2    : out    vl_logic;
        isEA_27DlyL2    : out    vl_logic;
        isEaMuxSel      : out    vl_logic;
        lcarE2          : out    vl_logic;
        lcarMuxSel      : out    vl_logic_vector(0 to 1);
        mux048Sel       : out    vl_logic_vector(0 to 1);
        nxtSwapSt       : out    vl_logic;
        pfb0BrTarSel    : out    vl_logic_vector(0 to 1);
        pfb0DataMuxSel  : out    vl_logic_vector(0 to 1);
        pfb0E1          : out    vl_logic;
        pfb0E2          : out    vl_logic;
        pfb0FullL2      : out    vl_logic;
        pfb0IarMuxSel   : out    vl_logic_vector(0 to 1);
        pfb1DataMuxSel  : out    vl_logic;
        pfb1E2          : out    vl_logic;
        pfb1IarMuxSel   : out    vl_logic;
        refetchAddrSel  : out    vl_logic;
        refetchLcarMuxSel: out    vl_logic_vector(0 to 1);
        refetchPipeStageSel: out    vl_logic_vector(0 to 1);
        runStL2         : out    vl_logic;
        saveForTraceE1  : out    vl_logic;
        saveForTraceE2  : out    vl_logic;
        seCtrSt         : out    vl_logic;
        seIdleSt        : out    vl_logic;
        stepStL2        : out    vl_logic;
        stuffStL2       : out    vl_logic;
        swapStL2        : out    vl_logic;
        traceDataSel    : out    vl_logic_vector(0 to 1);
        tracePipeHold   : out    vl_logic;
        tracePipeStageSel: out    vl_logic_vector(0 to 1);
        wbDataE1        : out    vl_logic;
        wbDataE2        : out    vl_logic;
        wbFlushOrClear  : out    vl_logic;
        wbIarE1         : out    vl_logic;
        wbIarE2         : out    vl_logic;
        APU_dcdValidOp_Neg: in     vl_logic;
        APU_sleepReq    : in     vl_logic;
        CB              : in     vl_logic;
        DBG_immdTE      : in     vl_logic_vector(0 to 2);
        DBG_stopReq     : in     vl_logic;
        DBG_wbTE        : in     vl_logic_vector(0 to 4);
        DBG_weakStopReq : in     vl_logic;
        DCU_sleepReq    : in     vl_logic;
        ICU_ifbE        : in     vl_logic;
        ICU_ifbO        : in     vl_logic;
        ICU_isCA        : in     vl_logic;
        ICU_sleepReq    : in     vl_logic;
        ICU_syncAfterReset: in     vl_logic;
        ICU_traceEnable : in     vl_logic;
        JTG_dbdrPulse   : in     vl_logic;
        JTG_step        : in     vl_logic;
        JTG_stopReq     : in     vl_logic;
        JTG_stuff       : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        MMU_isStatus    : in     vl_logic_vector(0 to 1);
        PCL_blkFlush    : in     vl_logic;
        PCL_dIcmpForStep: in     vl_logic;
        PCL_dIcmpForStuff: in     vl_logic;
        PCL_dcdHoldForIFB: in     vl_logic_vector(0 to 2);
        PCL_exe2Full    : in     vl_logic;
        PCL_exeIarHold  : in     vl_logic;
        PCL_icuOp_0     : in     vl_logic;
        PCL_wbClearTerms: in     vl_logic;
        PCL_wbFull      : in     vl_logic;
        PCL_wbHold      : in     vl_logic;
        PCL_wbStorageEnd: in     vl_logic;
        PCL_wbStorageOp : in     vl_logic;
        PGM_apuPresent  : in     vl_logic;
        TRC_fifoFull    : in     vl_logic;
        TRC_fifoOneEntryFree: in     vl_logic;
        TRC_se          : in     vl_logic;
        TRC_seCtrEqZeroL2: in     vl_logic;
        TRC_sleepReq    : in     vl_logic;
        VCT_anySwap     : in     vl_logic;
        VCT_msrWE       : in     vl_logic;
        VCT_swap01      : in     vl_logic;
        VCT_swap23      : in     vl_logic;
        VCT_wbFlush     : in     vl_logic;
        VCT_wbRfci      : in     vl_logic;
        VCT_wbRfi       : in     vl_logic;
        VCT_wbSuppress  : in     vl_logic;
        XXX_traceDisable: in     vl_logic;
        branchTarCrt    : in     vl_logic;
        coreReset       : in     vl_logic;
        dcdCorrect_Neg  : in     vl_logic;
        dcdData_5       : in     vl_logic;
        dcdData_21      : in     vl_logic;
        dcdData_30      : in     vl_logic;
        dcdTarget_Neg   : in     vl_logic;
        exeCorrect_Neg  : in     vl_logic;
        exeIsyncL2      : in     vl_logic;
        exeMtCtr        : in     vl_logic;
        exeMtLr         : in     vl_logic;
        exeRfciL2       : in     vl_logic;
        exeRfiL2        : in     vl_logic;
        exeScL2         : in     vl_logic;
        isEA_22         : in     vl_logic;
        isEA_27         : in     vl_logic;
        isEA_29         : in     vl_logic;
        lcar_29         : in     vl_logic;
        pfb0Data_5      : in     vl_logic;
        pfb0Data_21     : in     vl_logic;
        pfb0Data_30     : in     vl_logic;
        pfb0Target_Neg  : in     vl_logic;
        wbBrTakenL2     : in     vl_logic;
        wbIsyncL2       : in     vl_logic;
        wbMtCtrL2       : in     vl_logic;
        wbMtLrL2        : in     vl_logic;
        wbTEL2          : in     vl_logic_vector(0 to 4);
        MMU_isParityErr : in     vl_logic
    );
end p405s_fetcherCntl;
