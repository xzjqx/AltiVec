library verilog;
use verilog.vl_types.all;
entity p405s_exe_top is
    port(
        EXE_admMco      : out    vl_logic;
        EXE_apuLoadData : out    vl_logic_vector(0 to 31);
        EXE_cc          : out    vl_logic_vector(0 to 3);
        EXE_dac1CO      : out    vl_logic;
        EXE_dac1SumBit30Eq: out    vl_logic;
        EXE_dac1SumBit31Eq: out    vl_logic;
        EXE_dac1SumBits0thru27Eq: out    vl_logic;
        EXE_dac1SumBits28and29Eq: out    vl_logic;
        EXE_dac2CO      : out    vl_logic;
        EXE_dac2SumBit30Eq: out    vl_logic;
        EXE_dac2SumBit31Eq: out    vl_logic;
        EXE_dac2SumBits0thru27Eq: out    vl_logic;
        EXE_dac2SumBits28and29Eq: out    vl_logic;
        EXE_dcrAddr     : out    vl_logic_vector(0 to 9);
        EXE_dcrDataBus  : out    vl_logic_vector(0 to 31);
        EXE_dcuData     : out    vl_logic_vector(0 to 31);
        EXE_divMco      : out    vl_logic;
        EXE_dsEA_NEG    : out    vl_logic_vector(0 to 31);
        EXE_dsEaCP_NEG  : out    vl_logic_vector(0 to 7);
        EXE_dvc1ByteCmp : out    vl_logic_vector(0 to 3);
        EXE_dvc2ByteCmp : out    vl_logic_vector(0 to 3);
        EXE_ea          : out    vl_logic_vector(30 to 31);
        EXE_eaARegBuf   : out    vl_logic_vector(0 to 21);
        EXE_eaBRegBuf   : out    vl_logic_vector(0 to 21);
        EXE_ifbSprDataBus: out    vl_logic_vector(0 to 31);
        EXE_mmuIcuSprDataBus: out    vl_logic_vector(0 to 31);
        EXE_multMco     : out    vl_logic;
        EXE_raData      : out    vl_logic_vector(0 to 31);
        EXE_rbData      : out    vl_logic_vector(0 to 31);
        EXE_sprAddr     : out    vl_logic_vector(4 to 9);
        EXE_timJtgSprDataBus: out    vl_logic_vector(0 to 31);
        EXE_trap        : out    vl_logic;
        EXE_vctDbgSprDataBus: out    vl_logic_vector(0 to 31);
        EXE_wrteeIn     : out    vl_logic;
        EXE_xer         : out    vl_logic_vector(0 to 2);
        EXE_xerCa       : out    vl_logic;
        EXE_xerTBC      : out    vl_logic_vector(0 to 6);
        EXE_xerTBCIn    : out    vl_logic_vector(0 to 6);
        EXE_xerTBCNotEqZero: out    vl_logic;
        APU_exeCa       : in     vl_logic;
        APU_exeCr       : in     vl_logic_vector(0 to 3);
        APU_exeOv       : in     vl_logic;
        APU_exeResult   : in     vl_logic_vector(0 to 31);
        CB              : in     vl_logic;
        DBG_dacEn       : in     vl_logic;
        DBG_sprDataBus  : in     vl_logic_vector(0 to 31);
        DCU_SDQ_mod_NEG : in     vl_logic_vector(0 to 31);
        DCU_data_NEG    : in     vl_logic_vector(0 to 31);
        ICU_sprDataBus  : in     vl_logic_vector(0 to 31);
        IFB_exeMcrxr    : in     vl_logic;
        IFB_exeOpForExe2L2: in     vl_logic;
        IFB_sprDataBus  : in     vl_logic_vector(0 to 31);
        JTG_sprDataBus  : in     vl_logic_vector(0 to 31);
        LSSD_coreTestEn : in     vl_logic;
        MMU_sprDataBus  : in     vl_logic_vector(0 to 31);
        OCM_dsData      : in     vl_logic_vector(0 to 31);
        PCL_aPortRregBypass: in     vl_logic;
        PCL_aRegE2      : in     vl_logic;
        PCL_aRegForEaE2 : in     vl_logic;
        PCL_abRegE1     : in     vl_logic;
        PCL_addFour     : in     vl_logic;
        PCL_apuTrcLoadEn: in     vl_logic;
        PCL_bPortLitGenSel: in     vl_logic;
        PCL_bPortRregBypass: in     vl_logic;
        PCL_bRegE2      : in     vl_logic;
        PCL_bRegForEaE2 : in     vl_logic;
        PCL_dRegBypassMuxSel: in     vl_logic;
        PCL_dRegE1      : in     vl_logic;
        PCL_dbgSprDcds  : in     vl_logic_vector(0 to 3);
        PCL_dcdApAddr   : in     vl_logic_vector(0 to 9);
        PCL_dcdAregLoadUse: in     vl_logic;
        PCL_dcdBpAddr   : in     vl_logic_vector(0 to 9);
        PCL_dcdBregLoadUse: in     vl_logic;
        PCL_dcdHotCIn   : in     vl_logic;
        PCL_dcdImmd     : in     vl_logic_vector(11 to 31);
        PCL_dcdLitCntl  : in     vl_logic_vector(0 to 4);
        PCL_dcdMdSelQ   : in     vl_logic;
        PCL_dcdMrSelQ   : in     vl_logic;
        PCL_dcdSpAddr   : in     vl_logic_vector(0 to 9);
        PCL_dcdSregLoadUse: in     vl_logic;
        PCL_dcdSrmBpSel : in     vl_logic_vector(0 to 2);
        PCL_dcdXerCa    : in     vl_logic;
        PCL_dofDregE1   : in     vl_logic;
        PCL_dofDregMuxSel: in     vl_logic_vector(0 to 1);
        PCL_dvcByteEnL2 : in     vl_logic_vector(0 to 3);
        PCL_dvcCmpEn    : in     vl_logic;
        PCL_exe2AccRegMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exe2Hold    : in     vl_logic;
        PCL_exe2MacEn   : in     vl_logic;
        PCL_exe2MacOrMultEnForMS: in     vl_logic_vector(0 to 1);
        PCL_exe2MacOrMultEn_NEG: in     vl_logic_vector(0 to 1);
        PCL_exe2MacSat  : in     vl_logic;
        PCL_exe2MultEn  : in     vl_logic;
        PCL_exe2MultHiWd: in     vl_logic;
        PCL_exe2NegMac  : in     vl_logic;
        PCL_exe2SignedOp: in     vl_logic;
        PCL_exe2XerOvEn : in     vl_logic;
        PCL_exeAddEn    : in     vl_logic;
        PCL_exeAddSgndOp_NEG: in     vl_logic_vector(0 to 1);
        PCL_exeAdmCntl  : in     vl_logic_vector(0 to 3);
        PCL_exeApuValidOp: in     vl_logic;
        PCL_exeAregLoadUse: in     vl_logic;
        PCL_exeBregLoadUse: in     vl_logic;
        PCL_exeCmplmntA : in     vl_logic;
        PCL_exeCmplmntA_NEG: in     vl_logic;
        PCL_exeDivEn    : in     vl_logic;
        PCL_exeDivEnForLSSD: in     vl_logic;
        PCL_exeDivEnForMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exeDivEn_NEG: in     vl_logic;
        PCL_exeDivSgndOp: in     vl_logic;
        PCL_exeDvcHold  : in     vl_logic;
        PCL_exeEaCalc   : in     vl_logic;
        PCL_exeEaQwEn   : in     vl_logic_vector(0 to 3);
        PCL_exeFpuOp    : in     vl_logic;
        PCL_exeLoadUseHold: in     vl_logic;
        PCL_exeLogicalCntl: in     vl_logic_vector(0 to 7);
        PCL_exeLogicalUnitEnForLSSD: in     vl_logic;
        PCL_exeLogicalUnitEn_NEG: in     vl_logic;
        PCL_exeMacEn    : in     vl_logic;
        PCL_exeMacOrMultEn_NEG: in     vl_logic;
        PCL_exeMfspr    : in     vl_logic;
        PCL_exeMtspr    : in     vl_logic;
        PCL_exeMultEn   : in     vl_logic;
        PCL_exeMultEnForMuxSel: in     vl_logic_vector(0 to 1);
        PCL_exeMultEn_NEG: in     vl_logic_vector(0 to 1);
        PCL_exeNegMac   : in     vl_logic;
        PCL_exeRaEn     : in     vl_logic_vector(0 to 3);
        PCL_exeRbEn     : in     vl_logic_vector(0 to 3);
        PCL_exeSprDataEn_NEG: in     vl_logic;
        PCL_exeSprDcds  : in     vl_logic_vector(0 to 4);
        PCL_exeSprUnitEn_NEG: in     vl_logic;
        PCL_exeSregLoadUse: in     vl_logic;
        PCL_exeSrmBpSel : in     vl_logic_vector(0 to 2);
        PCL_exeSrmCntl  : in     vl_logic_vector(0 to 3);
        PCL_exeSrmUnitEnForLSSD: in     vl_logic;
        PCL_exeSrmUnitEn_NEG: in     vl_logic;
        PCL_exeTrapCond : in     vl_logic_vector(0 to 4);
        PCL_exeWrtee    : in     vl_logic;
        PCL_exeXerCaEn  : in     vl_logic;
        PCL_exeXerOvEn  : in     vl_logic;
        PCL_gateZeroToAreg: in     vl_logic;
        PCL_gateZeroToSreg: in     vl_logic;
        PCL_holdCIn     : in     vl_logic;
        PCL_holdMdMr    : in     vl_logic;
        PCL_ldAdjE1     : in     vl_logic;
        PCL_ldAdjE2     : in     vl_logic_vector(1 to 3);
        PCL_ldAdjMuxSel : in     vl_logic_vector(0 to 1);
        PCL_ldFillByPassMuxSel: in     vl_logic_vector(0 to 5);
        PCL_ldMuxSel    : in     vl_logic_vector(0 to 7);
        PCL_ldSteerMuxSel: in     vl_logic_vector(0 to 7);
        PCL_lwbLpAddr   : in     vl_logic_vector(0 to 4);
        PCL_lwbLpEqdcdApAddr: in     vl_logic;
        PCL_lwbLpEqdcdBpAddr: in     vl_logic;
        PCL_lwbLpEqdcdSpAddr: in     vl_logic;
        PCL_lwbLpWrEn   : in     vl_logic;
        PCL_mfDCRL2     : in     vl_logic;
        PCL_resultMuxSel: in     vl_logic;
        PCL_resultRegE1 : in     vl_logic;
        PCL_resultRegE2 : in     vl_logic;
        PCL_sPortRregBypass: in     vl_logic;
        PCL_sRegE1      : in     vl_logic;
        PCL_sRegE2      : in     vl_logic;
        PCL_sdqMuxSel   : in     vl_logic;
        PCL_sprHold     : in     vl_logic;
        PCL_sraRegE1    : in     vl_logic;
        PCL_sraRegE2    : in     vl_logic;
        PCL_srmRegE1    : in     vl_logic;
        PCL_srmRegE2    : in     vl_logic_vector(0 to 2);
        PCL_timSprDcds  : in     vl_logic_vector(0 to 5);
        PCL_vctSprDcds  : in     vl_logic_vector(0 to 5);
        PCL_wbHold      : in     vl_logic;
        PCL_wbRpAddr    : in     vl_logic_vector(0 to 4);
        PCL_wbRpEqdcdApAddr: in     vl_logic;
        PCL_wbRpEqdcdBpAddr: in     vl_logic;
        PCL_wbRpEqdcdSpAddr: in     vl_logic;
        PCL_wbRpWrEn    : in     vl_logic;
        PCL_xerL2Hold   : in     vl_logic;
        PGM_deterministicMult: in     vl_logic;
        TIM_sprDataBus  : in     vl_logic_vector(0 to 31);
        VCT_sprDataBus  : in     vl_logic_vector(0 to 31);
        XXX_dcrDataBus  : in     vl_logic_vector(0 to 31);
        coreReset       : in     vl_logic;
        PCL_exeDvcOrParityHold: in     vl_logic;
        DCU_parityError : in     vl_logic;
        EXE_dofDregParityErrL2: out    vl_logic;
        PCL_BpEqSp      : in     vl_logic;
        EXE_gprSysClkPI : in     vl_logic;
        EXE_gprRen      : in     vl_logic
    );
end p405s_exe_top;
