// 
// ************************************************************************** 
// 
//  Copyright (c) International Business Machines Corporation, 2005. 
// 
//  This file contains trade secrets and other proprietary and confidential 
//  information of International Business Machines Corporation which are 
//  protected by copyright and other intellectual property rights and shall 
//  not be reproduced, transferred to other documents, disclosed to others, 
//  or used for any purpose except as specifically authorized in writing by 
//  International Business Machines Corporation. This notice must be 
//  contained as part of this text at all times. 
// 
// ************************************************************************** 
//

module PPC405F5V1( C405APUDCDFULL, C405APUDCDHOLD, C405APUDCDINSTRUCTION00,
     C405APUDCDINSTRUCTION01, C405APUDCDINSTRUCTION02, C405APUDCDINSTRUCTION03,
     C405APUDCDINSTRUCTION04, C405APUDCDINSTRUCTION05, C405APUDCDINSTRUCTION06,
     C405APUDCDINSTRUCTION07, C405APUDCDINSTRUCTION08, C405APUDCDINSTRUCTION09,
     C405APUDCDINSTRUCTION10, C405APUDCDINSTRUCTION11, C405APUDCDINSTRUCTION12,
     C405APUDCDINSTRUCTION13, C405APUDCDINSTRUCTION14, C405APUDCDINSTRUCTION15,
     C405APUDCDINSTRUCTION16, C405APUDCDINSTRUCTION17, C405APUDCDINSTRUCTION18,
     C405APUDCDINSTRUCTION19, C405APUDCDINSTRUCTION20, C405APUDCDINSTRUCTION21,
     C405APUDCDINSTRUCTION22, C405APUDCDINSTRUCTION23, C405APUDCDINSTRUCTION24,
     C405APUDCDINSTRUCTION25, C405APUDCDINSTRUCTION26, C405APUDCDINSTRUCTION27,
     C405APUDCDINSTRUCTION28, C405APUDCDINSTRUCTION29, C405APUDCDINSTRUCTION30,
     C405APUDCDINSTRUCTION31, C405APUEXEFLUSH, C405APUEXEHOLD, C405APUEXELOADDBUS00,
     C405APUEXELOADDBUS01, C405APUEXELOADDBUS02, C405APUEXELOADDBUS03, C405APUEXELOADDBUS04,
     C405APUEXELOADDBUS05, C405APUEXELOADDBUS06, C405APUEXELOADDBUS07, C405APUEXELOADDBUS08,
     C405APUEXELOADDBUS09, C405APUEXELOADDBUS10, C405APUEXELOADDBUS11, C405APUEXELOADDBUS12,
     C405APUEXELOADDBUS13, C405APUEXELOADDBUS14, C405APUEXELOADDBUS15, C405APUEXELOADDBUS16,
     C405APUEXELOADDBUS17, C405APUEXELOADDBUS18, C405APUEXELOADDBUS19, C405APUEXELOADDBUS20,
     C405APUEXELOADDBUS21, C405APUEXELOADDBUS22, C405APUEXELOADDBUS23, C405APUEXELOADDBUS24,
     C405APUEXELOADDBUS25, C405APUEXELOADDBUS26, C405APUEXELOADDBUS27, C405APUEXELOADDBUS28,
     C405APUEXELOADDBUS29, C405APUEXELOADDBUS30, C405APUEXELOADDBUS31, C405APUEXELOADDVALID,
     C405APUEXERADATA00, C405APUEXERADATA01, C405APUEXERADATA02, C405APUEXERADATA03,
     C405APUEXERADATA04, C405APUEXERADATA05, C405APUEXERADATA06, C405APUEXERADATA07,
     C405APUEXERADATA08, C405APUEXERADATA09, C405APUEXERADATA10, C405APUEXERADATA11,
     C405APUEXERADATA12, C405APUEXERADATA13, C405APUEXERADATA14, C405APUEXERADATA15,
     C405APUEXERADATA16, C405APUEXERADATA17, C405APUEXERADATA18, C405APUEXERADATA19,
     C405APUEXERADATA20, C405APUEXERADATA21, C405APUEXERADATA22, C405APUEXERADATA23,
     C405APUEXERADATA24, C405APUEXERADATA25, C405APUEXERADATA26, C405APUEXERADATA27,
     C405APUEXERADATA28, C405APUEXERADATA29, C405APUEXERADATA30, C405APUEXERADATA31,
     C405APUEXERBDATA00, C405APUEXERBDATA01, C405APUEXERBDATA02, C405APUEXERBDATA03,
     C405APUEXERBDATA04, C405APUEXERBDATA05, C405APUEXERBDATA06, C405APUEXERBDATA07,
     C405APUEXERBDATA08, C405APUEXERBDATA09, C405APUEXERBDATA10, C405APUEXERBDATA11,
     C405APUEXERBDATA12, C405APUEXERBDATA13, C405APUEXERBDATA14, C405APUEXERBDATA15,
     C405APUEXERBDATA16, C405APUEXERBDATA17, C405APUEXERBDATA18, C405APUEXERBDATA19,
     C405APUEXERBDATA20, C405APUEXERBDATA21, C405APUEXERBDATA22, C405APUEXERBDATA23,
     C405APUEXERBDATA24, C405APUEXERBDATA25, C405APUEXERBDATA26, C405APUEXERBDATA27,
     C405APUEXERBDATA28, C405APUEXERBDATA29, C405APUEXERBDATA30, C405APUEXERBDATA31,
     C405APUEXEWDCNT0, C405APUEXEWDCNT1, C405APUMSRFE0, C405APUMSRFE1, C405APUWBBYTEEN0,
     C405APUWBBYTEEN1, C405APUWBBYTEEN2, C405APUWBBYTEEN3, C405APUWBENDIAN, C405APUWBFLUSH,
     C405APUWBHOLD, C405APUXERCA, C405CPMCORESLEEPREQ, C405CPMMSRCE, C405CPMMSREE,
     C405CPMTIMERIRQ, C405CPMTIMERRESETREQ, C405DBGLOADDATAONAPUDBUS, C405DBGMSRWE,
     C405DBGSTOPACK, C405DBGWBCOMPLETE, C405DBGWBFULL, C405DBGWBIAR00, C405DBGWBIAR01,
     C405DBGWBIAR02, C405DBGWBIAR03, C405DBGWBIAR04, C405DBGWBIAR05, C405DBGWBIAR06,
     C405DBGWBIAR07, C405DBGWBIAR08, C405DBGWBIAR09, C405DBGWBIAR10, C405DBGWBIAR11,
     C405DBGWBIAR12, C405DBGWBIAR13, C405DBGWBIAR14, C405DBGWBIAR15, C405DBGWBIAR16,
     C405DBGWBIAR17, C405DBGWBIAR18, C405DBGWBIAR19, C405DBGWBIAR20, C405DBGWBIAR21,
     C405DBGWBIAR22, C405DBGWBIAR23, C405DBGWBIAR24, C405DBGWBIAR25, C405DBGWBIAR26,
     C405DBGWBIAR27, C405DBGWBIAR28, C405DBGWBIAR29, C405DCRABUS0, C405DCRABUS1, C405DCRABUS2,
     C405DCRABUS3, C405DCRABUS4, C405DCRABUS5, C405DCRABUS6, C405DCRABUS7, C405DCRABUS8,
     C405DCRABUS9, C405DCRDBUSOUT00, C405DCRDBUSOUT01, C405DCRDBUSOUT02, C405DCRDBUSOUT03,
     C405DCRDBUSOUT04, C405DCRDBUSOUT05, C405DCRDBUSOUT06, C405DCRDBUSOUT07, C405DCRDBUSOUT08,
     C405DCRDBUSOUT09, C405DCRDBUSOUT10, C405DCRDBUSOUT11, C405DCRDBUSOUT12, C405DCRDBUSOUT13,
     C405DCRDBUSOUT14, C405DCRDBUSOUT15, C405DCRDBUSOUT16, C405DCRDBUSOUT17, C405DCRDBUSOUT18,
     C405DCRDBUSOUT19, C405DCRDBUSOUT20, C405DCRDBUSOUT21, C405DCRDBUSOUT22, C405DCRDBUSOUT23,
     C405DCRDBUSOUT24, C405DCRDBUSOUT25, C405DCRDBUSOUT26, C405DCRDBUSOUT27, C405DCRDBUSOUT28,
     C405DCRDBUSOUT29, C405DCRDBUSOUT30, C405DCRDBUSOUT31, C405DCRREAD, C405DCRWRITE,
     C405DSOCMABORTOP, C405DSOCMABORTREQ, C405DSOCMABUS00, C405DSOCMABUS01, C405DSOCMABUS02,
     C405DSOCMABUS03, C405DSOCMABUS04, C405DSOCMABUS05, C405DSOCMABUS06, C405DSOCMABUS07,
     C405DSOCMABUS08, C405DSOCMABUS09, C405DSOCMABUS10, C405DSOCMABUS11, C405DSOCMABUS12,
     C405DSOCMABUS13, C405DSOCMABUS14, C405DSOCMABUS15, C405DSOCMABUS16, C405DSOCMABUS17,
     C405DSOCMABUS18, C405DSOCMABUS19, C405DSOCMABUS20, C405DSOCMABUS21, C405DSOCMABUS22,
     C405DSOCMABUS23, C405DSOCMABUS24, C405DSOCMABUS25, C405DSOCMABUS26, C405DSOCMABUS27,
     C405DSOCMABUS28, C405DSOCMABUS29, C405DSOCMBYTEEN0, C405DSOCMBYTEEN1, C405DSOCMBYTEEN2,
     C405DSOCMBYTEEN3, C405DSOCMCACHEABLE, C405DSOCMGUARDED, C405DSOCMLOADREQ,
     C405DSOCMSTOREREQ, C405DSOCMSTRINGMULTIPLE, C405DSOCMU0ATTR, C405DSOCMWAIT,
     C405DSOCMWRDBUS00, C405DSOCMWRDBUS01, C405DSOCMWRDBUS02, C405DSOCMWRDBUS03,
     C405DSOCMWRDBUS04, C405DSOCMWRDBUS05, C405DSOCMWRDBUS06, C405DSOCMWRDBUS07,
     C405DSOCMWRDBUS08, C405DSOCMWRDBUS09, C405DSOCMWRDBUS10, C405DSOCMWRDBUS11,
     C405DSOCMWRDBUS12, C405DSOCMWRDBUS13, C405DSOCMWRDBUS14, C405DSOCMWRDBUS15,
     C405DSOCMWRDBUS16, C405DSOCMWRDBUS17, C405DSOCMWRDBUS18, C405DSOCMWRDBUS19,
     C405DSOCMWRDBUS20, C405DSOCMWRDBUS21, C405DSOCMWRDBUS22, C405DSOCMWRDBUS23,
     C405DSOCMWRDBUS24, C405DSOCMWRDBUS25, C405DSOCMWRDBUS26, C405DSOCMWRDBUS27,
     C405DSOCMWRDBUS28, C405DSOCMWRDBUS29, C405DSOCMWRDBUS30, C405DSOCMWRDBUS31,
     C405DSOCMXLATEVALID, C405ISOCMABORT, C405ISOCMABUS00, C405ISOCMABUS01, C405ISOCMABUS02,
     C405ISOCMABUS03, C405ISOCMABUS04, C405ISOCMABUS05, C405ISOCMABUS06, C405ISOCMABUS07,
     C405ISOCMABUS08, C405ISOCMABUS09, C405ISOCMABUS10, C405ISOCMABUS11, C405ISOCMABUS12,
     C405ISOCMABUS13, C405ISOCMABUS14, C405ISOCMABUS15, C405ISOCMABUS16, C405ISOCMABUS17,
     C405ISOCMABUS18, C405ISOCMABUS19, C405ISOCMABUS20, C405ISOCMABUS21, C405ISOCMABUS22,
     C405ISOCMABUS23, C405ISOCMABUS24, C405ISOCMABUS25, C405ISOCMABUS26, C405ISOCMABUS27,
     C405ISOCMABUS28, C405ISOCMABUS29, C405ISOCMCACHEABLE, C405ISOCMCONTEXTSYNC,
     C405ISOCMICUREADY, C405ISOCMREQPENDING, C405ISOCMU0ATTR, C405ISOCMXLATEVALID,
     C405JTGCAPTUREDR, C405JTGEXTEST, C405JTGPGMOUT, C405JTGSHIFTDR, C405JTGTDO, C405JTGTDOEN,
     C405JTGUPDATEDR, C405TESTDIAGABISTDONE,  C405TESTSCANOUT0,
     C405TESTSCANOUT1, C405TESTSCANOUT2, C405TESTSCANOUT3, C405TESTSCANOUT4, C405TESTSCANOUT5,
     C405TESTSCANOUT6, C405TESTSCANOUT7, C405PLBDCUABORT,
     C405PLBDCUABUS00, C405PLBDCUABUS01, C405PLBDCUABUS02, C405PLBDCUABUS03, C405PLBDCUABUS04,
     C405PLBDCUABUS05, C405PLBDCUABUS06, C405PLBDCUABUS07, C405PLBDCUABUS08, C405PLBDCUABUS09,
     C405PLBDCUABUS10, C405PLBDCUABUS11, C405PLBDCUABUS12, C405PLBDCUABUS13, C405PLBDCUABUS14,
     C405PLBDCUABUS15, C405PLBDCUABUS16, C405PLBDCUABUS17, C405PLBDCUABUS18, C405PLBDCUABUS19,
     C405PLBDCUABUS20, C405PLBDCUABUS21, C405PLBDCUABUS22, C405PLBDCUABUS23, C405PLBDCUABUS24,
     C405PLBDCUABUS25, C405PLBDCUABUS26, C405PLBDCUABUS27, C405PLBDCUABUS28, C405PLBDCUABUS29,
     C405PLBDCUABUS30, C405PLBDCUABUS31, C405PLBDCUBE0, C405PLBDCUBE1, C405PLBDCUBE2,
     C405PLBDCUBE3, C405PLBDCUBE4, C405PLBDCUBE5, C405PLBDCUBE6, C405PLBDCUBE7,
     C405PLBDCUCACHEABLE, C405PLBDCUGUARDED, C405PLBDCUPRIORITY0, C405PLBDCUPRIORITY1,
     C405PLBDCUREQUEST, C405PLBDCURNW, C405PLBDCUSIZE2, C405PLBDCUU0ATTR, C405PLBDCUWRDBUS00,
     C405PLBDCUWRDBUS01, C405PLBDCUWRDBUS02, C405PLBDCUWRDBUS03, C405PLBDCUWRDBUS04,
     C405PLBDCUWRDBUS05, C405PLBDCUWRDBUS06, C405PLBDCUWRDBUS07, C405PLBDCUWRDBUS08,
     C405PLBDCUWRDBUS09, C405PLBDCUWRDBUS10, C405PLBDCUWRDBUS11, C405PLBDCUWRDBUS12,
     C405PLBDCUWRDBUS13, C405PLBDCUWRDBUS14, C405PLBDCUWRDBUS15, C405PLBDCUWRDBUS16,
     C405PLBDCUWRDBUS17, C405PLBDCUWRDBUS18, C405PLBDCUWRDBUS19, C405PLBDCUWRDBUS20,
     C405PLBDCUWRDBUS21, C405PLBDCUWRDBUS22, C405PLBDCUWRDBUS23, C405PLBDCUWRDBUS24,
     C405PLBDCUWRDBUS25, C405PLBDCUWRDBUS26, C405PLBDCUWRDBUS27, C405PLBDCUWRDBUS28,
     C405PLBDCUWRDBUS29, C405PLBDCUWRDBUS30, C405PLBDCUWRDBUS31, C405PLBDCUWRDBUS32,
     C405PLBDCUWRDBUS33, C405PLBDCUWRDBUS34, C405PLBDCUWRDBUS35, C405PLBDCUWRDBUS36,
     C405PLBDCUWRDBUS37, C405PLBDCUWRDBUS38, C405PLBDCUWRDBUS39, C405PLBDCUWRDBUS40,
     C405PLBDCUWRDBUS41, C405PLBDCUWRDBUS42, C405PLBDCUWRDBUS43, C405PLBDCUWRDBUS44,
     C405PLBDCUWRDBUS45, C405PLBDCUWRDBUS46, C405PLBDCUWRDBUS47, C405PLBDCUWRDBUS48,
     C405PLBDCUWRDBUS49, C405PLBDCUWRDBUS50, C405PLBDCUWRDBUS51, C405PLBDCUWRDBUS52,
     C405PLBDCUWRDBUS53, C405PLBDCUWRDBUS54, C405PLBDCUWRDBUS55, C405PLBDCUWRDBUS56,
     C405PLBDCUWRDBUS57, C405PLBDCUWRDBUS58, C405PLBDCUWRDBUS59, C405PLBDCUWRDBUS60,
     C405PLBDCUWRDBUS61, C405PLBDCUWRDBUS62, C405PLBDCUWRDBUS63, C405PLBDCUWRITETHRU,
     C405PLBICUABORT, C405PLBICUABUS00, C405PLBICUABUS01, C405PLBICUABUS02, C405PLBICUABUS03,
     C405PLBICUABUS04, C405PLBICUABUS05, C405PLBICUABUS06, C405PLBICUABUS07, C405PLBICUABUS08,
     C405PLBICUABUS09, C405PLBICUABUS10, C405PLBICUABUS11, C405PLBICUABUS12, C405PLBICUABUS13,
     C405PLBICUABUS14, C405PLBICUABUS15, C405PLBICUABUS16, C405PLBICUABUS17, C405PLBICUABUS18,
     C405PLBICUABUS19, C405PLBICUABUS20, C405PLBICUABUS21, C405PLBICUABUS22, C405PLBICUABUS23,
     C405PLBICUABUS24, C405PLBICUABUS25, C405PLBICUABUS26, C405PLBICUABUS27, C405PLBICUABUS28,
     C405PLBICUABUS29, C405PLBICUCACHEABLE, C405PLBICUPRIORITY0, C405PLBICUPRIORITY1,
     C405PLBICUREQUEST, C405PLBICUSIZE2, C405PLBICUSIZE3, C405PLBICUU0ATTR,
     C405RSTCHIPRESETREQ, C405RSTCORERESETREQ, C405RSTSYSTEMRESETREQ, C405TRCCYCLE,
     C405TRCEVENEXECUTIONSTATUS0, C405TRCEVENEXECUTIONSTATUS1, C405TRCODDEXECUTIONSTATUS0,
     C405TRCODDEXECUTIONSTATUS1, C405TRCTRACESTATUS0, C405TRCTRACESTATUS1, C405TRCTRACESTATUS2,
     C405TRCTRACESTATUS3, C405TRCTRIGGEREVENTOUT, C405TRCTRIGGEREVENTTYPE0,
     C405TRCTRIGGEREVENTTYPE1, C405TRCTRIGGEREVENTTYPE2, C405TRCTRIGGEREVENTTYPE3,
     C405TRCTRIGGEREVENTTYPE4, C405TRCTRIGGEREVENTTYPE5, C405TRCTRIGGEREVENTTYPE6,
     C405TRCTRIGGEREVENTTYPE7, C405TRCTRIGGEREVENTTYPE8, C405TRCTRIGGEREVENTTYPE9,
     C405TRCTRIGGEREVENTTYPE10, C405XXXMACHINECHECK, APUC405DCDAPUOP, APUC405DCDCREN,
     APUC405DCDFORCEALGN, APUC405DCDFORCEBESTEERING, APUC405DCDFPUOP, APUC405DCDGPRWRITE,
     APUC405DCDLDSTBYTE, APUC405DCDLDSTDW, APUC405DCDLDSTHW, APUC405DCDLDSTQW,
     APUC405DCDLDSTWD, APUC405DCDLOAD, APUC405DCDPRIVOP, APUC405DCDRAEN, APUC405DCDRBEN,
     APUC405DCDSTORE, APUC405DCDTRAPBE, APUC405DCDTRAPLE, APUC405DCDUPDATE, APUC405DCDVALIDOP,
     APUC405DCDXERCAEN, APUC405DCDXEROVEN, APUC405EXCEPTION, APUC405EXEBLOCKINGMCO,
     APUC405EXEBUSY, APUC405EXECR0, APUC405EXECR1, APUC405EXECR2, APUC405EXECR3,
     APUC405EXECRFIELD0, APUC405EXECRFIELD1, APUC405EXECRFIELD2, APUC405EXELDDEPEND,
     APUC405EXENONBLOCKINGMCO, APUC405EXERESULT00, APUC405EXERESULT01, APUC405EXERESULT02,
     APUC405EXERESULT03, APUC405EXERESULT04, APUC405EXERESULT05, APUC405EXERESULT06,
     APUC405EXERESULT07, APUC405EXERESULT08, APUC405EXERESULT09, APUC405EXERESULT10,
     APUC405EXERESULT11, APUC405EXERESULT12, APUC405EXERESULT13, APUC405EXERESULT14,
     APUC405EXERESULT15, APUC405EXERESULT16, APUC405EXERESULT17, APUC405EXERESULT18,
     APUC405EXERESULT19, APUC405EXERESULT20, APUC405EXERESULT21, APUC405EXERESULT22,
     APUC405EXERESULT23, APUC405EXERESULT24, APUC405EXERESULT25, APUC405EXERESULT26,
     APUC405EXERESULT27, APUC405EXERESULT28, APUC405EXERESULT29, APUC405EXERESULT30,
     APUC405EXERESULT31, APUC405EXEXERCA, APUC405EXEXEROV, APUC405FPUEXCEPTION,
     APUC405LWBLDDEPEND, APUC405SLEEPREQ, APUC405WBLDDEPEND, CPMC405CLOCK, CPMC405CPUCLKENCCLK,
     CPMC405CORECLKINACTIVE,  CPMC405JTAGCLKENCCLK,
     CPMC405PLBSAMPLECYCLE, CPMC405TIMERCLKENCCLK, CPMC405TIMERTICK, DBGC405DEBUGHALT,
     DBGC405EXTBUSHOLDACK, DBGC405UNCONDDEBUGEVENT, DCRC405ACK, DCRC405DBUSIN00,
     DCRC405DBUSIN01, DCRC405DBUSIN02, DCRC405DBUSIN03, DCRC405DBUSIN04, DCRC405DBUSIN05,
     DCRC405DBUSIN06, DCRC405DBUSIN07, DCRC405DBUSIN08, DCRC405DBUSIN09, DCRC405DBUSIN10,
     DCRC405DBUSIN11, DCRC405DBUSIN12, DCRC405DBUSIN13, DCRC405DBUSIN14, DCRC405DBUSIN15,
     DCRC405DBUSIN16, DCRC405DBUSIN17, DCRC405DBUSIN18, DCRC405DBUSIN19, DCRC405DBUSIN20,
     DCRC405DBUSIN21, DCRC405DBUSIN22, DCRC405DBUSIN23, DCRC405DBUSIN24, DCRC405DBUSIN25,
     DCRC405DBUSIN26, DCRC405DBUSIN27, DCRC405DBUSIN28, DCRC405DBUSIN29, DCRC405DBUSIN30,
     DCRC405DBUSIN31, DSOCMC405COMPLETE, DSOCMC405DISOPERANDFWD, DSOCMC405HOLD,
     DSOCMC405RDDBUS00, DSOCMC405RDDBUS01, DSOCMC405RDDBUS02, DSOCMC405RDDBUS03,
     DSOCMC405RDDBUS04, DSOCMC405RDDBUS05, DSOCMC405RDDBUS06, DSOCMC405RDDBUS07,
     DSOCMC405RDDBUS08, DSOCMC405RDDBUS09, DSOCMC405RDDBUS10, DSOCMC405RDDBUS11,
     DSOCMC405RDDBUS12, DSOCMC405RDDBUS13, DSOCMC405RDDBUS14, DSOCMC405RDDBUS15,
     DSOCMC405RDDBUS16, DSOCMC405RDDBUS17, DSOCMC405RDDBUS18, DSOCMC405RDDBUS19,
     DSOCMC405RDDBUS20, DSOCMC405RDDBUS21, DSOCMC405RDDBUS22, DSOCMC405RDDBUS23,
     DSOCMC405RDDBUS24, DSOCMC405RDDBUS25, DSOCMC405RDDBUS26, DSOCMC405RDDBUS27,
     DSOCMC405RDDBUS28, DSOCMC405RDDBUS29, DSOCMC405RDDBUS30, DSOCMC405RDDBUS31,
     EICC405CRITINPUTIRQ, EICC405EXTINPUTIRQ, ISOCMC405HOLD, ISOCMC405RDDBUS00,
     ISOCMC405RDDBUS01, ISOCMC405RDDBUS02, ISOCMC405RDDBUS03, ISOCMC405RDDBUS04,
     ISOCMC405RDDBUS05, ISOCMC405RDDBUS06, ISOCMC405RDDBUS07, ISOCMC405RDDBUS08,
     ISOCMC405RDDBUS09, ISOCMC405RDDBUS10, ISOCMC405RDDBUS11, ISOCMC405RDDBUS12,
     ISOCMC405RDDBUS13, ISOCMC405RDDBUS14, ISOCMC405RDDBUS15, ISOCMC405RDDBUS16,
     ISOCMC405RDDBUS17, ISOCMC405RDDBUS18, ISOCMC405RDDBUS19, ISOCMC405RDDBUS20,
     ISOCMC405RDDBUS21, ISOCMC405RDDBUS22, ISOCMC405RDDBUS23, ISOCMC405RDDBUS24,
     ISOCMC405RDDBUS25, ISOCMC405RDDBUS26, ISOCMC405RDDBUS27, ISOCMC405RDDBUS28,
     ISOCMC405RDDBUS29, ISOCMC405RDDBUS30, ISOCMC405RDDBUS31, ISOCMC405RDDBUS32,
     ISOCMC405RDDBUS33, ISOCMC405RDDBUS34, ISOCMC405RDDBUS35, ISOCMC405RDDBUS36,
     ISOCMC405RDDBUS37, ISOCMC405RDDBUS38, ISOCMC405RDDBUS39, ISOCMC405RDDBUS40,
     ISOCMC405RDDBUS41, ISOCMC405RDDBUS42, ISOCMC405RDDBUS43, ISOCMC405RDDBUS44,
     ISOCMC405RDDBUS45, ISOCMC405RDDBUS46, ISOCMC405RDDBUS47, ISOCMC405RDDBUS48,
     ISOCMC405RDDBUS49, ISOCMC405RDDBUS50, ISOCMC405RDDBUS51, ISOCMC405RDDBUS52,
     ISOCMC405RDDBUS53, ISOCMC405RDDBUS54, ISOCMC405RDDBUS55, ISOCMC405RDDBUS56,
     ISOCMC405RDDBUS57, ISOCMC405RDDBUS58, ISOCMC405RDDBUS59, ISOCMC405RDDBUS60,
     ISOCMC405RDDBUS61, ISOCMC405RDDBUS62, ISOCMC405RDDBUS63, ISOCMC405RDDVALID0,
     ISOCMC405RDDVALID1, JTGC405BNDSCANTDO, JTGC405TCK, JTGC405TDI, JTGC405TMS, JTGC405TRSTNEG,
     TESTC405BISTCCLK, 
     TESTC405SCANIN0, TESTC405SCANIN1, TESTC405SCANIN2, TESTC405SCANIN3, TESTC405SCANIN4,
     TESTC405SCANIN5, TESTC405SCANIN6, TESTC405SCANIN7, TESTC405SCANENABLE, TESTC405TESTMODE,
     TESTC405CNTLPOINT, TESTC405TESTM1, TESTC405TESTM3, PLBC405DCUADDRACK, PLBC405DCUBUSY,
     PLBC405DCUERR, PLBC405DCURDDACK, PLBC405DCURDDBUS00, PLBC405DCURDDBUS01,
     PLBC405DCURDDBUS02, PLBC405DCURDDBUS03, PLBC405DCURDDBUS04, PLBC405DCURDDBUS05,
     PLBC405DCURDDBUS06, PLBC405DCURDDBUS07, PLBC405DCURDDBUS08, PLBC405DCURDDBUS09,
     PLBC405DCURDDBUS10, PLBC405DCURDDBUS11, PLBC405DCURDDBUS12, PLBC405DCURDDBUS13,
     PLBC405DCURDDBUS14, PLBC405DCURDDBUS15, PLBC405DCURDDBUS16, PLBC405DCURDDBUS17,
     PLBC405DCURDDBUS18, PLBC405DCURDDBUS19, PLBC405DCURDDBUS20, PLBC405DCURDDBUS21,
     PLBC405DCURDDBUS22, PLBC405DCURDDBUS23, PLBC405DCURDDBUS24, PLBC405DCURDDBUS25,
     PLBC405DCURDDBUS26, PLBC405DCURDDBUS27, PLBC405DCURDDBUS28, PLBC405DCURDDBUS29,
     PLBC405DCURDDBUS30, PLBC405DCURDDBUS31, PLBC405DCURDDBUS32, PLBC405DCURDDBUS33,
     PLBC405DCURDDBUS34, PLBC405DCURDDBUS35, PLBC405DCURDDBUS36, PLBC405DCURDDBUS37,
     PLBC405DCURDDBUS38, PLBC405DCURDDBUS39, PLBC405DCURDDBUS40, PLBC405DCURDDBUS41,
     PLBC405DCURDDBUS42, PLBC405DCURDDBUS43, PLBC405DCURDDBUS44, PLBC405DCURDDBUS45,
     PLBC405DCURDDBUS46, PLBC405DCURDDBUS47, PLBC405DCURDDBUS48, PLBC405DCURDDBUS49,
     PLBC405DCURDDBUS50, PLBC405DCURDDBUS51, PLBC405DCURDDBUS52, PLBC405DCURDDBUS53,
     PLBC405DCURDDBUS54, PLBC405DCURDDBUS55, PLBC405DCURDDBUS56, PLBC405DCURDDBUS57,
     PLBC405DCURDDBUS58, PLBC405DCURDDBUS59, PLBC405DCURDDBUS60, PLBC405DCURDDBUS61,
     PLBC405DCURDDBUS62, PLBC405DCURDDBUS63, PLBC405DCURDWDADDR1, PLBC405DCURDWDADDR2,
     PLBC405DCURDWDADDR3, PLBC405DCUSSIZE1, PLBC405DCUWRDACK, PLBC405ICUADDRACK,
     PLBC405ICUBUSY, PLBC405ICUERR, PLBC405ICURDDACK, PLBC405ICURDDBUS00, PLBC405ICURDDBUS01,
     PLBC405ICURDDBUS02, PLBC405ICURDDBUS03, PLBC405ICURDDBUS04, PLBC405ICURDDBUS05,
     PLBC405ICURDDBUS06, PLBC405ICURDDBUS07, PLBC405ICURDDBUS08, PLBC405ICURDDBUS09,
     PLBC405ICURDDBUS10, PLBC405ICURDDBUS11, PLBC405ICURDDBUS12, PLBC405ICURDDBUS13,
     PLBC405ICURDDBUS14, PLBC405ICURDDBUS15, PLBC405ICURDDBUS16, PLBC405ICURDDBUS17,
     PLBC405ICURDDBUS18, PLBC405ICURDDBUS19, PLBC405ICURDDBUS20, PLBC405ICURDDBUS21,
     PLBC405ICURDDBUS22, PLBC405ICURDDBUS23, PLBC405ICURDDBUS24, PLBC405ICURDDBUS25,
     PLBC405ICURDDBUS26, PLBC405ICURDDBUS27, PLBC405ICURDDBUS28, PLBC405ICURDDBUS29,
     PLBC405ICURDDBUS30, PLBC405ICURDDBUS31, PLBC405ICURDDBUS32, PLBC405ICURDDBUS33,
     PLBC405ICURDDBUS34, PLBC405ICURDDBUS35, PLBC405ICURDDBUS36, PLBC405ICURDDBUS37,
     PLBC405ICURDDBUS38, PLBC405ICURDDBUS39, PLBC405ICURDDBUS40, PLBC405ICURDDBUS41,
     PLBC405ICURDDBUS42, PLBC405ICURDDBUS43, PLBC405ICURDDBUS44, PLBC405ICURDDBUS45,
     PLBC405ICURDDBUS46, PLBC405ICURDDBUS47, PLBC405ICURDDBUS48, PLBC405ICURDDBUS49,
     PLBC405ICURDDBUS50, PLBC405ICURDDBUS51, PLBC405ICURDDBUS52, PLBC405ICURDDBUS53,
     PLBC405ICURDDBUS54, PLBC405ICURDDBUS55, PLBC405ICURDDBUS56, PLBC405ICURDDBUS57,
     PLBC405ICURDDBUS58, PLBC405ICURDDBUS59, PLBC405ICURDDBUS60, PLBC405ICURDDBUS61,
     PLBC405ICURDDBUS62, PLBC405ICURDDBUS63, PLBC405ICURDWDADDR1, PLBC405ICURDWDADDR2,
     PLBC405ICURDWDADDR3, PLBC405ICUSSIZE1, RSTC405RESETCHIP, RSTC405RESETCORE,
     RSTC405RESETSYSTEM, TIEC405APUDIVEN, TIEC405APUPRESENT, TIEC405DETERMINISTICMULT,
     TIEC405DISOPERANDFWD, TIEC405MMUEN, TIEC405PVR00, TIEC405PVR01, TIEC405PVR02,
     TIEC405PVR03, TIEC405PVR04, TIEC405PVR05, TIEC405PVR06, TIEC405PVR07, TIEC405PVR08,
     TIEC405PVR09, TIEC405PVR10, TIEC405PVR11, TIEC405PVR12, TIEC405PVR13, TIEC405PVR14,
     TIEC405PVR15, TIEC405PVR16, TIEC405PVR17, TIEC405PVR18, TIEC405PVR19, TIEC405PVR20,
     TIEC405PVR21, TIEC405PVR22, TIEC405PVR23, TIEC405PVR24, TIEC405PVR25, TIEC405PVR26,
     TIEC405PVR27, TIEC405PVR28, TIEC405PVR29, TIEC405PVR30, TIEC405PVR31, TRCC405TRACEDISABLE,
     TRCC405TRIGGEREVENTIN, 
     C405BISTPEPSPF00, C405BISTPEPSPF01,
     C405BISTPEPSPF02, TESTC405CE0EVS, TESTC405BISTCE0STCLK,
     TESTC405BISTCE1ENABLE,  TESTC405BISTCE1MODE, 
     CPMC405PLBSYNCCLOCK, CPMC405SYNCBYPASS, TIEC405CLOCKENABLE, TIEC405DUTYENABLE,
     CPMC405PLBSAMPLECYCLEALT,
     BISTC405DCUBISTDEBUGSI00,BISTC405DCUBISTDEBUGSI01, BISTC405DCUBISTDEBUGSI02, BISTC405DCUBISTDEBUGSI03,
     C405BISTDCUBISTDEBUGSO00, C405BISTDCUBISTDEBUGSO01,C405BISTDCUBISTDEBUGSO02,C405BISTDCUBISTDEBUGSO03,
     BISTC405DCUBISTDEBUGEN00,BISTC405DCUBISTDEBUGEN01,BISTC405DCUBISTDEBUGEN02,BISTC405DCUBISTDEBUGEN03,
     BISTC405DCUBISTMODEREGIN00,BISTC405DCUBISTMODEREGIN01,BISTC405DCUBISTMODEREGIN02,
     BISTC405DCUBISTMODEREGIN03,BISTC405DCUBISTMODEREGIN04,BISTC405DCUBISTMODEREGIN05,
     BISTC405DCUBISTMODEREGIN06,BISTC405DCUBISTMODEREGIN07,BISTC405DCUBISTMODEREGIN08,
     BISTC405DCUBISTMODEREGIN09,BISTC405DCUBISTMODEREGIN10,BISTC405DCUBISTMODEREGIN11,
     BISTC405DCUBISTMODEREGIN12,BISTC405DCUBISTMODEREGIN13,BISTC405DCUBISTMODEREGIN14,
     BISTC405DCUBISTMODEREGIN15,BISTC405DCUBISTMODEREGIN16,BISTC405DCUBISTMODEREGIN17,
     BISTC405DCUBISTMODEREGIN18,
     C405BISTDCUBISTMODEREGOUT00,C405BISTDCUBISTMODEREGOUT01,C405BISTDCUBISTMODEREGOUT02,
     C405BISTDCUBISTMODEREGOUT03,C405BISTDCUBISTMODEREGOUT04,C405BISTDCUBISTMODEREGOUT05,
     C405BISTDCUBISTMODEREGOUT06,C405BISTDCUBISTMODEREGOUT07,C405BISTDCUBISTMODEREGOUT08,
     C405BISTDCUBISTMODEREGOUT09,C405BISTDCUBISTMODEREGOUT10,C405BISTDCUBISTMODEREGOUT11,
     C405BISTDCUBISTMODEREGOUT12,C405BISTDCUBISTMODEREGOUT13,C405BISTDCUBISTMODEREGOUT14,
     C405BISTDCUBISTMODEREGOUT15,C405BISTDCUBISTMODEREGOUT16,C405BISTDCUBISTMODEREGOUT17,
     C405BISTDCUBISTMODEREGOUT18,
     BISTC405DCUBISTMODEREGSI,
     C405BISTDCUBISTMODEREGSO,
     BISTC405DCUBISTSHIFTDR,
     BISTC405DCUBISTMBRUN,
     BISTC405DCUBISTPARALLELDR,

     BISTC405ICUBISTDEBUGSI00,BISTC405ICUBISTDEBUGSI01, BISTC405ICUBISTDEBUGSI02, BISTC405ICUBISTDEBUGSI03,
     C405BISTICUBISTDEBUGSO00, C405BISTICUBISTDEBUGSO01,C405BISTICUBISTDEBUGSO02,C405BISTICUBISTDEBUGSO03,
     BISTC405ICUBISTDEBUGEN00,BISTC405ICUBISTDEBUGEN01,BISTC405ICUBISTDEBUGEN02,BISTC405ICUBISTDEBUGEN03,
     BISTC405ICUBISTMODEREGIN00,BISTC405ICUBISTMODEREGIN01,BISTC405ICUBISTMODEREGIN02,
     BISTC405ICUBISTMODEREGIN03,BISTC405ICUBISTMODEREGIN04,BISTC405ICUBISTMODEREGIN05,
     BISTC405ICUBISTMODEREGIN06,BISTC405ICUBISTMODEREGIN07,BISTC405ICUBISTMODEREGIN08,
     BISTC405ICUBISTMODEREGIN09,BISTC405ICUBISTMODEREGIN10,BISTC405ICUBISTMODEREGIN11,
     BISTC405ICUBISTMODEREGIN12,BISTC405ICUBISTMODEREGIN13,BISTC405ICUBISTMODEREGIN14,
     BISTC405ICUBISTMODEREGIN15,BISTC405ICUBISTMODEREGIN16,BISTC405ICUBISTMODEREGIN17,
     BISTC405ICUBISTMODEREGIN18,
     C405BISTICUBISTMODEREGOUT00,C405BISTICUBISTMODEREGOUT01,C405BISTICUBISTMODEREGOUT02,
     C405BISTICUBISTMODEREGOUT03,C405BISTICUBISTMODEREGOUT04,C405BISTICUBISTMODEREGOUT05,
     C405BISTICUBISTMODEREGOUT06,C405BISTICUBISTMODEREGOUT07,C405BISTICUBISTMODEREGOUT08,
     C405BISTICUBISTMODEREGOUT09,C405BISTICUBISTMODEREGOUT10,C405BISTICUBISTMODEREGOUT11,
     C405BISTICUBISTMODEREGOUT12,C405BISTICUBISTMODEREGOUT13,C405BISTICUBISTMODEREGOUT14,
     C405BISTICUBISTMODEREGOUT15,C405BISTICUBISTMODEREGOUT16,C405BISTICUBISTMODEREGOUT17,
     C405BISTICUBISTMODEREGOUT18,
     BISTC405ICUBISTMODEREGSI,
     C405BISTICUBISTMODEREGSO,
     BISTC405ICUBISTSHIFTDR,
     BISTC405ICUBISTMBRUN,
     BISTC405ICUBISTPARALLELDR
   );
     
output  C405APUDCDFULL, C405APUDCDHOLD, C405APUDCDINSTRUCTION00, C405APUDCDINSTRUCTION01,
     C405APUDCDINSTRUCTION02, C405APUDCDINSTRUCTION03, C405APUDCDINSTRUCTION04,
     C405APUDCDINSTRUCTION05, C405APUDCDINSTRUCTION06, C405APUDCDINSTRUCTION07,
     C405APUDCDINSTRUCTION08, C405APUDCDINSTRUCTION09, C405APUDCDINSTRUCTION10,
     C405APUDCDINSTRUCTION11, C405APUDCDINSTRUCTION12, C405APUDCDINSTRUCTION13,
     C405APUDCDINSTRUCTION14, C405APUDCDINSTRUCTION15, C405APUDCDINSTRUCTION16,
     C405APUDCDINSTRUCTION17, C405APUDCDINSTRUCTION18, C405APUDCDINSTRUCTION19,
     C405APUDCDINSTRUCTION20, C405APUDCDINSTRUCTION21, C405APUDCDINSTRUCTION22,
     C405APUDCDINSTRUCTION23, C405APUDCDINSTRUCTION24, C405APUDCDINSTRUCTION25,
     C405APUDCDINSTRUCTION26, C405APUDCDINSTRUCTION27, C405APUDCDINSTRUCTION28,
     C405APUDCDINSTRUCTION29, C405APUDCDINSTRUCTION30, C405APUDCDINSTRUCTION31,
     C405APUEXEFLUSH, C405APUEXEHOLD, C405APUEXELOADDBUS00, C405APUEXELOADDBUS01,
     C405APUEXELOADDBUS02, C405APUEXELOADDBUS03, C405APUEXELOADDBUS04, C405APUEXELOADDBUS05,
     C405APUEXELOADDBUS06, C405APUEXELOADDBUS07, C405APUEXELOADDBUS08, C405APUEXELOADDBUS09,
     C405APUEXELOADDBUS10, C405APUEXELOADDBUS11, C405APUEXELOADDBUS12, C405APUEXELOADDBUS13,
     C405APUEXELOADDBUS14, C405APUEXELOADDBUS15, C405APUEXELOADDBUS16, C405APUEXELOADDBUS17,
     C405APUEXELOADDBUS18, C405APUEXELOADDBUS19, C405APUEXELOADDBUS20, C405APUEXELOADDBUS21,
     C405APUEXELOADDBUS22, C405APUEXELOADDBUS23, C405APUEXELOADDBUS24, C405APUEXELOADDBUS25,
     C405APUEXELOADDBUS26, C405APUEXELOADDBUS27, C405APUEXELOADDBUS28, C405APUEXELOADDBUS29,
     C405APUEXELOADDBUS30, C405APUEXELOADDBUS31, C405APUEXELOADDVALID, C405APUEXERADATA00,
     C405APUEXERADATA01, C405APUEXERADATA02, C405APUEXERADATA03, C405APUEXERADATA04,
     C405APUEXERADATA05, C405APUEXERADATA06, C405APUEXERADATA07, C405APUEXERADATA08,
     C405APUEXERADATA09, C405APUEXERADATA10, C405APUEXERADATA11, C405APUEXERADATA12,
     C405APUEXERADATA13, C405APUEXERADATA14, C405APUEXERADATA15, C405APUEXERADATA16,
     C405APUEXERADATA17, C405APUEXERADATA18, C405APUEXERADATA19, C405APUEXERADATA20,
     C405APUEXERADATA21, C405APUEXERADATA22, C405APUEXERADATA23, C405APUEXERADATA24,
     C405APUEXERADATA25, C405APUEXERADATA26, C405APUEXERADATA27, C405APUEXERADATA28,
     C405APUEXERADATA29, C405APUEXERADATA30, C405APUEXERADATA31, C405APUEXERBDATA00,
     C405APUEXERBDATA01, C405APUEXERBDATA02, C405APUEXERBDATA03, C405APUEXERBDATA04,
     C405APUEXERBDATA05, C405APUEXERBDATA06, C405APUEXERBDATA07, C405APUEXERBDATA08,
     C405APUEXERBDATA09, C405APUEXERBDATA10, C405APUEXERBDATA11, C405APUEXERBDATA12,
     C405APUEXERBDATA13, C405APUEXERBDATA14, C405APUEXERBDATA15, C405APUEXERBDATA16,
     C405APUEXERBDATA17, C405APUEXERBDATA18, C405APUEXERBDATA19, C405APUEXERBDATA20,
     C405APUEXERBDATA21, C405APUEXERBDATA22, C405APUEXERBDATA23, C405APUEXERBDATA24,
     C405APUEXERBDATA25, C405APUEXERBDATA26, C405APUEXERBDATA27, C405APUEXERBDATA28,
     C405APUEXERBDATA29, C405APUEXERBDATA30, C405APUEXERBDATA31, C405APUEXEWDCNT0,
     C405APUEXEWDCNT1, C405APUMSRFE0, C405APUMSRFE1, C405APUWBBYTEEN0, C405APUWBBYTEEN1,
     C405APUWBBYTEEN2, C405APUWBBYTEEN3, C405APUWBENDIAN, C405APUWBFLUSH, C405APUWBHOLD,
     C405APUXERCA, C405CPMCORESLEEPREQ, C405CPMMSRCE, C405CPMMSREE, C405CPMTIMERIRQ,
     C405CPMTIMERRESETREQ, C405DBGLOADDATAONAPUDBUS, C405DBGMSRWE, C405DBGSTOPACK,
     C405DBGWBCOMPLETE, C405DBGWBFULL, C405DBGWBIAR00, C405DBGWBIAR01, C405DBGWBIAR02,
     C405DBGWBIAR03, C405DBGWBIAR04, C405DBGWBIAR05, C405DBGWBIAR06, C405DBGWBIAR07,
     C405DBGWBIAR08, C405DBGWBIAR09, C405DBGWBIAR10, C405DBGWBIAR11, C405DBGWBIAR12,
     C405DBGWBIAR13, C405DBGWBIAR14, C405DBGWBIAR15, C405DBGWBIAR16, C405DBGWBIAR17,
     C405DBGWBIAR18, C405DBGWBIAR19, C405DBGWBIAR20, C405DBGWBIAR21, C405DBGWBIAR22,
     C405DBGWBIAR23, C405DBGWBIAR24, C405DBGWBIAR25, C405DBGWBIAR26, C405DBGWBIAR27,
     C405DBGWBIAR28, C405DBGWBIAR29, C405DCRABUS0, C405DCRABUS1, C405DCRABUS2, C405DCRABUS3,
     C405DCRABUS4, C405DCRABUS5, C405DCRABUS6, C405DCRABUS7, C405DCRABUS8, C405DCRABUS9,
     C405DCRDBUSOUT00, C405DCRDBUSOUT01, C405DCRDBUSOUT02, C405DCRDBUSOUT03, C405DCRDBUSOUT04,
     C405DCRDBUSOUT05, C405DCRDBUSOUT06, C405DCRDBUSOUT07, C405DCRDBUSOUT08, C405DCRDBUSOUT09,
     C405DCRDBUSOUT10, C405DCRDBUSOUT11, C405DCRDBUSOUT12, C405DCRDBUSOUT13, C405DCRDBUSOUT14,
     C405DCRDBUSOUT15, C405DCRDBUSOUT16, C405DCRDBUSOUT17, C405DCRDBUSOUT18, C405DCRDBUSOUT19,
     C405DCRDBUSOUT20, C405DCRDBUSOUT21, C405DCRDBUSOUT22, C405DCRDBUSOUT23, C405DCRDBUSOUT24,
     C405DCRDBUSOUT25, C405DCRDBUSOUT26, C405DCRDBUSOUT27, C405DCRDBUSOUT28, C405DCRDBUSOUT29,
     C405DCRDBUSOUT30, C405DCRDBUSOUT31, C405DCRREAD, C405DCRWRITE, C405DSOCMABORTOP,
     C405DSOCMABORTREQ, C405DSOCMABUS00, C405DSOCMABUS01, C405DSOCMABUS02, C405DSOCMABUS03,
     C405DSOCMABUS04, C405DSOCMABUS05, C405DSOCMABUS06, C405DSOCMABUS07, C405DSOCMABUS08,
     C405DSOCMABUS09, C405DSOCMABUS10, C405DSOCMABUS11, C405DSOCMABUS12, C405DSOCMABUS13,
     C405DSOCMABUS14, C405DSOCMABUS15, C405DSOCMABUS16, C405DSOCMABUS17, C405DSOCMABUS18,
     C405DSOCMABUS19, C405DSOCMABUS20, C405DSOCMABUS21, C405DSOCMABUS22, C405DSOCMABUS23,
     C405DSOCMABUS24, C405DSOCMABUS25, C405DSOCMABUS26, C405DSOCMABUS27, C405DSOCMABUS28,
     C405DSOCMABUS29, C405DSOCMBYTEEN0, C405DSOCMBYTEEN1, C405DSOCMBYTEEN2, C405DSOCMBYTEEN3,
     C405DSOCMCACHEABLE, C405DSOCMGUARDED, C405DSOCMLOADREQ, C405DSOCMSTOREREQ,
     C405DSOCMSTRINGMULTIPLE, C405DSOCMU0ATTR, C405DSOCMWAIT, C405DSOCMWRDBUS00,
     C405DSOCMWRDBUS01, C405DSOCMWRDBUS02, C405DSOCMWRDBUS03, C405DSOCMWRDBUS04,
     C405DSOCMWRDBUS05, C405DSOCMWRDBUS06, C405DSOCMWRDBUS07, C405DSOCMWRDBUS08,
     C405DSOCMWRDBUS09, C405DSOCMWRDBUS10, C405DSOCMWRDBUS11, C405DSOCMWRDBUS12,
     C405DSOCMWRDBUS13, C405DSOCMWRDBUS14, C405DSOCMWRDBUS15, C405DSOCMWRDBUS16,
     C405DSOCMWRDBUS17, C405DSOCMWRDBUS18, C405DSOCMWRDBUS19, C405DSOCMWRDBUS20,
     C405DSOCMWRDBUS21, C405DSOCMWRDBUS22, C405DSOCMWRDBUS23, C405DSOCMWRDBUS24,
     C405DSOCMWRDBUS25, C405DSOCMWRDBUS26, C405DSOCMWRDBUS27, C405DSOCMWRDBUS28,
     C405DSOCMWRDBUS29, C405DSOCMWRDBUS30, C405DSOCMWRDBUS31, C405DSOCMXLATEVALID,
     C405ISOCMABORT, C405ISOCMABUS00, C405ISOCMABUS01, C405ISOCMABUS02, C405ISOCMABUS03,
     C405ISOCMABUS04, C405ISOCMABUS05, C405ISOCMABUS06, C405ISOCMABUS07, C405ISOCMABUS08,
     C405ISOCMABUS09, C405ISOCMABUS10, C405ISOCMABUS11, C405ISOCMABUS12, C405ISOCMABUS13,
     C405ISOCMABUS14, C405ISOCMABUS15, C405ISOCMABUS16, C405ISOCMABUS17, C405ISOCMABUS18,
     C405ISOCMABUS19, C405ISOCMABUS20, C405ISOCMABUS21, C405ISOCMABUS22, C405ISOCMABUS23,
     C405ISOCMABUS24, C405ISOCMABUS25, C405ISOCMABUS26, C405ISOCMABUS27, C405ISOCMABUS28,
     C405ISOCMABUS29, C405ISOCMCACHEABLE, C405ISOCMCONTEXTSYNC, C405ISOCMICUREADY,
     C405ISOCMREQPENDING, C405ISOCMU0ATTR, C405ISOCMXLATEVALID, C405JTGCAPTUREDR,
     C405JTGEXTEST, C405JTGPGMOUT, C405JTGSHIFTDR, C405JTGTDO, C405JTGTDOEN, C405JTGUPDATEDR,
     C405TESTDIAGABISTDONE,  C405TESTSCANOUT0, C405TESTSCANOUT1,
     C405TESTSCANOUT2, C405TESTSCANOUT3, C405TESTSCANOUT4, C405TESTSCANOUT5, C405TESTSCANOUT6,
     C405TESTSCANOUT7, C405PLBDCUABORT, C405PLBDCUABUS00,
     C405PLBDCUABUS01, C405PLBDCUABUS02, C405PLBDCUABUS03, C405PLBDCUABUS04, C405PLBDCUABUS05,
     C405PLBDCUABUS06, C405PLBDCUABUS07, C405PLBDCUABUS08, C405PLBDCUABUS09, C405PLBDCUABUS10,
     C405PLBDCUABUS11, C405PLBDCUABUS12, C405PLBDCUABUS13, C405PLBDCUABUS14, C405PLBDCUABUS15,
     C405PLBDCUABUS16, C405PLBDCUABUS17, C405PLBDCUABUS18, C405PLBDCUABUS19, C405PLBDCUABUS20,
     C405PLBDCUABUS21, C405PLBDCUABUS22, C405PLBDCUABUS23, C405PLBDCUABUS24, C405PLBDCUABUS25,
     C405PLBDCUABUS26, C405PLBDCUABUS27, C405PLBDCUABUS28, C405PLBDCUABUS29, C405PLBDCUABUS30,
     C405PLBDCUABUS31, C405PLBDCUBE0, C405PLBDCUBE1, C405PLBDCUBE2, C405PLBDCUBE3,
     C405PLBDCUBE4, C405PLBDCUBE5, C405PLBDCUBE6, C405PLBDCUBE7, C405PLBDCUCACHEABLE,
     C405PLBDCUGUARDED, C405PLBDCUPRIORITY0, C405PLBDCUPRIORITY1, C405PLBDCUREQUEST,
     C405PLBDCURNW, C405PLBDCUSIZE2, C405PLBDCUU0ATTR, C405PLBDCUWRDBUS00, C405PLBDCUWRDBUS01,
     C405PLBDCUWRDBUS02, C405PLBDCUWRDBUS03, C405PLBDCUWRDBUS04, C405PLBDCUWRDBUS05,
     C405PLBDCUWRDBUS06, C405PLBDCUWRDBUS07, C405PLBDCUWRDBUS08, C405PLBDCUWRDBUS09,
     C405PLBDCUWRDBUS10, C405PLBDCUWRDBUS11, C405PLBDCUWRDBUS12, C405PLBDCUWRDBUS13,
     C405PLBDCUWRDBUS14, C405PLBDCUWRDBUS15, C405PLBDCUWRDBUS16, C405PLBDCUWRDBUS17,
     C405PLBDCUWRDBUS18, C405PLBDCUWRDBUS19, C405PLBDCUWRDBUS20, C405PLBDCUWRDBUS21,
     C405PLBDCUWRDBUS22, C405PLBDCUWRDBUS23, C405PLBDCUWRDBUS24, C405PLBDCUWRDBUS25,
     C405PLBDCUWRDBUS26, C405PLBDCUWRDBUS27, C405PLBDCUWRDBUS28, C405PLBDCUWRDBUS29,
     C405PLBDCUWRDBUS30, C405PLBDCUWRDBUS31, C405PLBDCUWRDBUS32, C405PLBDCUWRDBUS33,
     C405PLBDCUWRDBUS34, C405PLBDCUWRDBUS35, C405PLBDCUWRDBUS36, C405PLBDCUWRDBUS37,
     C405PLBDCUWRDBUS38, C405PLBDCUWRDBUS39, C405PLBDCUWRDBUS40, C405PLBDCUWRDBUS41,
     C405PLBDCUWRDBUS42, C405PLBDCUWRDBUS43, C405PLBDCUWRDBUS44, C405PLBDCUWRDBUS45,
     C405PLBDCUWRDBUS46, C405PLBDCUWRDBUS47, C405PLBDCUWRDBUS48, C405PLBDCUWRDBUS49,
     C405PLBDCUWRDBUS50, C405PLBDCUWRDBUS51, C405PLBDCUWRDBUS52, C405PLBDCUWRDBUS53,
     C405PLBDCUWRDBUS54, C405PLBDCUWRDBUS55, C405PLBDCUWRDBUS56, C405PLBDCUWRDBUS57,
     C405PLBDCUWRDBUS58, C405PLBDCUWRDBUS59, C405PLBDCUWRDBUS60, C405PLBDCUWRDBUS61,
     C405PLBDCUWRDBUS62, C405PLBDCUWRDBUS63, C405PLBDCUWRITETHRU, C405PLBICUABORT,
     C405PLBICUABUS00, C405PLBICUABUS01, C405PLBICUABUS02, C405PLBICUABUS03, C405PLBICUABUS04,
     C405PLBICUABUS05, C405PLBICUABUS06, C405PLBICUABUS07, C405PLBICUABUS08, C405PLBICUABUS09,
     C405PLBICUABUS10, C405PLBICUABUS11, C405PLBICUABUS12, C405PLBICUABUS13, C405PLBICUABUS14,
     C405PLBICUABUS15, C405PLBICUABUS16, C405PLBICUABUS17, C405PLBICUABUS18, C405PLBICUABUS19,
     C405PLBICUABUS20, C405PLBICUABUS21, C405PLBICUABUS22, C405PLBICUABUS23, C405PLBICUABUS24,
     C405PLBICUABUS25, C405PLBICUABUS26, C405PLBICUABUS27, C405PLBICUABUS28, C405PLBICUABUS29,
     C405PLBICUCACHEABLE, C405PLBICUPRIORITY0, C405PLBICUPRIORITY1, C405PLBICUREQUEST,
     C405PLBICUSIZE2, C405PLBICUSIZE3, C405PLBICUU0ATTR, C405RSTCHIPRESETREQ,
     C405RSTCORERESETREQ, C405RSTSYSTEMRESETREQ, C405TRCCYCLE, C405TRCEVENEXECUTIONSTATUS0,
     C405TRCEVENEXECUTIONSTATUS1, C405TRCODDEXECUTIONSTATUS0, C405TRCODDEXECUTIONSTATUS1,
     C405TRCTRACESTATUS0, C405TRCTRACESTATUS1, C405TRCTRACESTATUS2, C405TRCTRACESTATUS3,
     C405TRCTRIGGEREVENTOUT, C405TRCTRIGGEREVENTTYPE0, C405TRCTRIGGEREVENTTYPE1,
     C405TRCTRIGGEREVENTTYPE2, C405TRCTRIGGEREVENTTYPE3, C405TRCTRIGGEREVENTTYPE4,
     C405TRCTRIGGEREVENTTYPE5, C405TRCTRIGGEREVENTTYPE6, C405TRCTRIGGEREVENTTYPE7,
     C405TRCTRIGGEREVENTTYPE8, C405TRCTRIGGEREVENTTYPE9, C405TRCTRIGGEREVENTTYPE10,
     C405XXXMACHINECHECK, 
     C405BISTPEPSPF00, C405BISTPEPSPF01, C405BISTPEPSPF02;


input  APUC405DCDAPUOP, APUC405DCDCREN, APUC405DCDFORCEALGN, APUC405DCDFORCEBESTEERING,
     APUC405DCDFPUOP, APUC405DCDGPRWRITE, APUC405DCDLDSTBYTE, APUC405DCDLDSTDW,
     APUC405DCDLDSTHW, APUC405DCDLDSTQW, APUC405DCDLDSTWD, APUC405DCDLOAD, APUC405DCDPRIVOP,
     APUC405DCDRAEN, APUC405DCDRBEN, APUC405DCDSTORE, APUC405DCDTRAPBE, APUC405DCDTRAPLE,
     APUC405DCDUPDATE, APUC405DCDVALIDOP, APUC405DCDXERCAEN, APUC405DCDXEROVEN,
     APUC405EXCEPTION, APUC405EXEBLOCKINGMCO, APUC405EXEBUSY, APUC405EXECR0, APUC405EXECR1,
     APUC405EXECR2, APUC405EXECR3, APUC405EXECRFIELD0, APUC405EXECRFIELD1, APUC405EXECRFIELD2,
     APUC405EXELDDEPEND, APUC405EXENONBLOCKINGMCO, APUC405EXERESULT00, APUC405EXERESULT01,
     APUC405EXERESULT02, APUC405EXERESULT03, APUC405EXERESULT04, APUC405EXERESULT05,
     APUC405EXERESULT06, APUC405EXERESULT07, APUC405EXERESULT08, APUC405EXERESULT09,
     APUC405EXERESULT10, APUC405EXERESULT11, APUC405EXERESULT12, APUC405EXERESULT13,
     APUC405EXERESULT14, APUC405EXERESULT15, APUC405EXERESULT16, APUC405EXERESULT17,
     APUC405EXERESULT18, APUC405EXERESULT19, APUC405EXERESULT20, APUC405EXERESULT21,
     APUC405EXERESULT22, APUC405EXERESULT23, APUC405EXERESULT24, APUC405EXERESULT25,
     APUC405EXERESULT26, APUC405EXERESULT27, APUC405EXERESULT28, APUC405EXERESULT29,
     APUC405EXERESULT30, APUC405EXERESULT31, APUC405EXEXERCA, APUC405EXEXEROV,
     APUC405FPUEXCEPTION, APUC405LWBLDDEPEND, APUC405SLEEPREQ, APUC405WBLDDEPEND, CPMC405CLOCK,
     CPMC405CPUCLKENCCLK, CPMC405CORECLKINACTIVE,  CPMC405JTAGCLKENCCLK,
     CPMC405PLBSAMPLECYCLE, CPMC405TIMERCLKENCCLK, CPMC405TIMERTICK, DBGC405DEBUGHALT,
     DBGC405EXTBUSHOLDACK, DBGC405UNCONDDEBUGEVENT, DCRC405ACK, DCRC405DBUSIN00,
     DCRC405DBUSIN01, DCRC405DBUSIN02, DCRC405DBUSIN03, DCRC405DBUSIN04, DCRC405DBUSIN05,
     DCRC405DBUSIN06, DCRC405DBUSIN07, DCRC405DBUSIN08, DCRC405DBUSIN09, DCRC405DBUSIN10,
     DCRC405DBUSIN11, DCRC405DBUSIN12, DCRC405DBUSIN13, DCRC405DBUSIN14, DCRC405DBUSIN15,
     DCRC405DBUSIN16, DCRC405DBUSIN17, DCRC405DBUSIN18, DCRC405DBUSIN19, DCRC405DBUSIN20,
     DCRC405DBUSIN21, DCRC405DBUSIN22, DCRC405DBUSIN23, DCRC405DBUSIN24, DCRC405DBUSIN25,
     DCRC405DBUSIN26, DCRC405DBUSIN27, DCRC405DBUSIN28, DCRC405DBUSIN29, DCRC405DBUSIN30,
     DCRC405DBUSIN31, DSOCMC405COMPLETE, DSOCMC405DISOPERANDFWD, DSOCMC405HOLD,
     DSOCMC405RDDBUS00, DSOCMC405RDDBUS01, DSOCMC405RDDBUS02, DSOCMC405RDDBUS03,
     DSOCMC405RDDBUS04, DSOCMC405RDDBUS05, DSOCMC405RDDBUS06, DSOCMC405RDDBUS07,
     DSOCMC405RDDBUS08, DSOCMC405RDDBUS09, DSOCMC405RDDBUS10, DSOCMC405RDDBUS11,
     DSOCMC405RDDBUS12, DSOCMC405RDDBUS13, DSOCMC405RDDBUS14, DSOCMC405RDDBUS15,
     DSOCMC405RDDBUS16, DSOCMC405RDDBUS17, DSOCMC405RDDBUS18, DSOCMC405RDDBUS19,
     DSOCMC405RDDBUS20, DSOCMC405RDDBUS21, DSOCMC405RDDBUS22, DSOCMC405RDDBUS23,
     DSOCMC405RDDBUS24, DSOCMC405RDDBUS25, DSOCMC405RDDBUS26, DSOCMC405RDDBUS27,
     DSOCMC405RDDBUS28, DSOCMC405RDDBUS29, DSOCMC405RDDBUS30, DSOCMC405RDDBUS31,
     EICC405CRITINPUTIRQ, EICC405EXTINPUTIRQ, ISOCMC405HOLD, ISOCMC405RDDBUS00,
     ISOCMC405RDDBUS01, ISOCMC405RDDBUS02, ISOCMC405RDDBUS03, ISOCMC405RDDBUS04,
     ISOCMC405RDDBUS05, ISOCMC405RDDBUS06, ISOCMC405RDDBUS07, ISOCMC405RDDBUS08,
     ISOCMC405RDDBUS09, ISOCMC405RDDBUS10, ISOCMC405RDDBUS11, ISOCMC405RDDBUS12,
     ISOCMC405RDDBUS13, ISOCMC405RDDBUS14, ISOCMC405RDDBUS15, ISOCMC405RDDBUS16,
     ISOCMC405RDDBUS17, ISOCMC405RDDBUS18, ISOCMC405RDDBUS19, ISOCMC405RDDBUS20,
     ISOCMC405RDDBUS21, ISOCMC405RDDBUS22, ISOCMC405RDDBUS23, ISOCMC405RDDBUS24,
     ISOCMC405RDDBUS25, ISOCMC405RDDBUS26, ISOCMC405RDDBUS27, ISOCMC405RDDBUS28,
     ISOCMC405RDDBUS29, ISOCMC405RDDBUS30, ISOCMC405RDDBUS31, ISOCMC405RDDBUS32,
     ISOCMC405RDDBUS33, ISOCMC405RDDBUS34, ISOCMC405RDDBUS35, ISOCMC405RDDBUS36,
     ISOCMC405RDDBUS37, ISOCMC405RDDBUS38, ISOCMC405RDDBUS39, ISOCMC405RDDBUS40,
     ISOCMC405RDDBUS41, ISOCMC405RDDBUS42, ISOCMC405RDDBUS43, ISOCMC405RDDBUS44,
     ISOCMC405RDDBUS45, ISOCMC405RDDBUS46, ISOCMC405RDDBUS47, ISOCMC405RDDBUS48,
     ISOCMC405RDDBUS49, ISOCMC405RDDBUS50, ISOCMC405RDDBUS51, ISOCMC405RDDBUS52,
     ISOCMC405RDDBUS53, ISOCMC405RDDBUS54, ISOCMC405RDDBUS55, ISOCMC405RDDBUS56,
     ISOCMC405RDDBUS57, ISOCMC405RDDBUS58, ISOCMC405RDDBUS59, ISOCMC405RDDBUS60,
     ISOCMC405RDDBUS61, ISOCMC405RDDBUS62, ISOCMC405RDDBUS63, ISOCMC405RDDVALID0,
     ISOCMC405RDDVALID1, JTGC405BNDSCANTDO, JTGC405TCK, JTGC405TDI, JTGC405TMS, JTGC405TRSTNEG,
     TESTC405BISTCCLK, 
     TESTC405SCANIN0, TESTC405SCANIN1, TESTC405SCANIN2, TESTC405SCANIN3, TESTC405SCANIN4,
     TESTC405SCANIN5, TESTC405SCANIN6, TESTC405SCANIN7, TESTC405SCANENABLE, TESTC405TESTMODE,
     TESTC405CNTLPOINT, TESTC405TESTM1, TESTC405TESTM3, PLBC405DCUADDRACK, PLBC405DCUBUSY,
     PLBC405DCUERR, PLBC405DCURDDACK, PLBC405DCURDDBUS00, PLBC405DCURDDBUS01,
     PLBC405DCURDDBUS02, PLBC405DCURDDBUS03, PLBC405DCURDDBUS04, PLBC405DCURDDBUS05,
     PLBC405DCURDDBUS06, PLBC405DCURDDBUS07, PLBC405DCURDDBUS08, PLBC405DCURDDBUS09,
     PLBC405DCURDDBUS10, PLBC405DCURDDBUS11, PLBC405DCURDDBUS12, PLBC405DCURDDBUS13,
     PLBC405DCURDDBUS14, PLBC405DCURDDBUS15, PLBC405DCURDDBUS16, PLBC405DCURDDBUS17,
     PLBC405DCURDDBUS18, PLBC405DCURDDBUS19, PLBC405DCURDDBUS20, PLBC405DCURDDBUS21,
     PLBC405DCURDDBUS22, PLBC405DCURDDBUS23, PLBC405DCURDDBUS24, PLBC405DCURDDBUS25,
     PLBC405DCURDDBUS26, PLBC405DCURDDBUS27, PLBC405DCURDDBUS28, PLBC405DCURDDBUS29,
     PLBC405DCURDDBUS30, PLBC405DCURDDBUS31, PLBC405DCURDDBUS32, PLBC405DCURDDBUS33,
     PLBC405DCURDDBUS34, PLBC405DCURDDBUS35, PLBC405DCURDDBUS36, PLBC405DCURDDBUS37,
     PLBC405DCURDDBUS38, PLBC405DCURDDBUS39, PLBC405DCURDDBUS40, PLBC405DCURDDBUS41,
     PLBC405DCURDDBUS42, PLBC405DCURDDBUS43, PLBC405DCURDDBUS44, PLBC405DCURDDBUS45,
     PLBC405DCURDDBUS46, PLBC405DCURDDBUS47, PLBC405DCURDDBUS48, PLBC405DCURDDBUS49,
     PLBC405DCURDDBUS50, PLBC405DCURDDBUS51, PLBC405DCURDDBUS52, PLBC405DCURDDBUS53,
     PLBC405DCURDDBUS54, PLBC405DCURDDBUS55, PLBC405DCURDDBUS56, PLBC405DCURDDBUS57,
     PLBC405DCURDDBUS58, PLBC405DCURDDBUS59, PLBC405DCURDDBUS60, PLBC405DCURDDBUS61,
     PLBC405DCURDDBUS62, PLBC405DCURDDBUS63, PLBC405DCURDWDADDR1, PLBC405DCURDWDADDR2,
     PLBC405DCURDWDADDR3, PLBC405DCUSSIZE1, PLBC405DCUWRDACK, PLBC405ICUADDRACK,
     PLBC405ICUBUSY, PLBC405ICUERR, PLBC405ICURDDACK, PLBC405ICURDDBUS00, PLBC405ICURDDBUS01,
     PLBC405ICURDDBUS02, PLBC405ICURDDBUS03, PLBC405ICURDDBUS04, PLBC405ICURDDBUS05,
     PLBC405ICURDDBUS06, PLBC405ICURDDBUS07, PLBC405ICURDDBUS08, PLBC405ICURDDBUS09,
     PLBC405ICURDDBUS10, PLBC405ICURDDBUS11, PLBC405ICURDDBUS12, PLBC405ICURDDBUS13,
     PLBC405ICURDDBUS14, PLBC405ICURDDBUS15, PLBC405ICURDDBUS16, PLBC405ICURDDBUS17,
     PLBC405ICURDDBUS18, PLBC405ICURDDBUS19, PLBC405ICURDDBUS20, PLBC405ICURDDBUS21,
     PLBC405ICURDDBUS22, PLBC405ICURDDBUS23, PLBC405ICURDDBUS24, PLBC405ICURDDBUS25,
     PLBC405ICURDDBUS26, PLBC405ICURDDBUS27, PLBC405ICURDDBUS28, PLBC405ICURDDBUS29,
     PLBC405ICURDDBUS30, PLBC405ICURDDBUS31, PLBC405ICURDDBUS32, PLBC405ICURDDBUS33,
     PLBC405ICURDDBUS34, PLBC405ICURDDBUS35, PLBC405ICURDDBUS36, PLBC405ICURDDBUS37,
     PLBC405ICURDDBUS38, PLBC405ICURDDBUS39, PLBC405ICURDDBUS40, PLBC405ICURDDBUS41,
     PLBC405ICURDDBUS42, PLBC405ICURDDBUS43, PLBC405ICURDDBUS44, PLBC405ICURDDBUS45,
     PLBC405ICURDDBUS46, PLBC405ICURDDBUS47, PLBC405ICURDDBUS48, PLBC405ICURDDBUS49,
     PLBC405ICURDDBUS50, PLBC405ICURDDBUS51, PLBC405ICURDDBUS52, PLBC405ICURDDBUS53,
     PLBC405ICURDDBUS54, PLBC405ICURDDBUS55, PLBC405ICURDDBUS56, PLBC405ICURDDBUS57,
     PLBC405ICURDDBUS58, PLBC405ICURDDBUS59, PLBC405ICURDDBUS60, PLBC405ICURDDBUS61,
     PLBC405ICURDDBUS62, PLBC405ICURDDBUS63, PLBC405ICURDWDADDR1, PLBC405ICURDWDADDR2,
     PLBC405ICURDWDADDR3, PLBC405ICUSSIZE1, RSTC405RESETCHIP, RSTC405RESETCORE,
     RSTC405RESETSYSTEM, TIEC405APUDIVEN, TIEC405APUPRESENT, TIEC405DETERMINISTICMULT,
     TIEC405DISOPERANDFWD, TIEC405MMUEN, TIEC405PVR00, TIEC405PVR01, TIEC405PVR02,
     TIEC405PVR03, TIEC405PVR04, TIEC405PVR05, TIEC405PVR06, TIEC405PVR07, TIEC405PVR08,
     TIEC405PVR09, TIEC405PVR10, TIEC405PVR11, TIEC405PVR12, TIEC405PVR13, TIEC405PVR14,
     TIEC405PVR15, TIEC405PVR16, TIEC405PVR17, TIEC405PVR18, TIEC405PVR19, TIEC405PVR20,
     TIEC405PVR21, TIEC405PVR22, TIEC405PVR23, TIEC405PVR24, TIEC405PVR25, TIEC405PVR26,
     TIEC405PVR27, TIEC405PVR28, TIEC405PVR29, TIEC405PVR30, TIEC405PVR31, TRCC405TRACEDISABLE,
     TRCC405TRIGGEREVENTIN, TESTC405CE0EVS, TESTC405BISTCE0STCLK,
     TESTC405BISTCE1ENABLE, TESTC405BISTCE1MODE, 
     CPMC405PLBSYNCCLOCK, CPMC405SYNCBYPASS, TIEC405CLOCKENABLE, TIEC405DUTYENABLE,
     CPMC405PLBSAMPLECYCLEALT;

// BIST Interface

input          BISTC405DCUBISTMBRUN;

//input  [3:0]   BISTC405DCUBISTDEBUGSI;
wire  [3:0]   dcu_bist_debug_si;
input     BISTC405DCUBISTDEBUGSI00;
input     BISTC405DCUBISTDEBUGSI01;
input     BISTC405DCUBISTDEBUGSI02;
input     BISTC405DCUBISTDEBUGSI03;
assign dcu_bist_debug_si = {BISTC405DCUBISTDEBUGSI00, BISTC405DCUBISTDEBUGSI01,BISTC405DCUBISTDEBUGSI02,BISTC405DCUBISTDEBUGSI03}; 
//input  [3:0]   BISTC405DCUBISTDEBUGEN;
wire  [3:0]   dcu_bist_debug_en;
input    BISTC405DCUBISTDEBUGEN00;
input    BISTC405DCUBISTDEBUGEN01;
input    BISTC405DCUBISTDEBUGEN02;
input    BISTC405DCUBISTDEBUGEN03;
assign dcu_bist_debug_en = { BISTC405DCUBISTDEBUGEN00, BISTC405DCUBISTDEBUGEN01, BISTC405DCUBISTDEBUGEN02, BISTC405DCUBISTDEBUGEN03};
//output [3:0]   C405BISTDCUBISTDEBUGSO;
wire [3:0]   dcu_bist_debug_so;
output   C405BISTDCUBISTDEBUGSO00;
output   C405BISTDCUBISTDEBUGSO01;
output   C405BISTDCUBISTDEBUGSO02;
output   C405BISTDCUBISTDEBUGSO03;
assign  {C405BISTDCUBISTDEBUGSO00, C405BISTDCUBISTDEBUGSO01,C405BISTDCUBISTDEBUGSO02,C405BISTDCUBISTDEBUGSO03} = dcu_bist_debug_so ;

input          BISTC405DCUBISTSHIFTDR;
input          BISTC405DCUBISTMODEREGSI;
output         C405BISTDCUBISTMODEREGSO;

input          BISTC405DCUBISTPARALLELDR;
input     BISTC405DCUBISTMODEREGIN00,BISTC405DCUBISTMODEREGIN01,BISTC405DCUBISTMODEREGIN02,
     BISTC405DCUBISTMODEREGIN03,BISTC405DCUBISTMODEREGIN04,BISTC405DCUBISTMODEREGIN05,
     BISTC405DCUBISTMODEREGIN06,BISTC405DCUBISTMODEREGIN07,BISTC405DCUBISTMODEREGIN08,
     BISTC405DCUBISTMODEREGIN09,BISTC405DCUBISTMODEREGIN10,BISTC405DCUBISTMODEREGIN11,
     BISTC405DCUBISTMODEREGIN12,BISTC405DCUBISTMODEREGIN13,BISTC405DCUBISTMODEREGIN14,
     BISTC405DCUBISTMODEREGIN15,BISTC405DCUBISTMODEREGIN16,BISTC405DCUBISTMODEREGIN17,
     BISTC405DCUBISTMODEREGIN18;
wire  [18:0]  dcu_bist_mode_reg_in;
assign dcu_bist_mode_reg_in = {
     BISTC405DCUBISTMODEREGIN00,BISTC405DCUBISTMODEREGIN01,BISTC405DCUBISTMODEREGIN02,
     BISTC405DCUBISTMODEREGIN03,BISTC405DCUBISTMODEREGIN04,BISTC405DCUBISTMODEREGIN05,
     BISTC405DCUBISTMODEREGIN06,BISTC405DCUBISTMODEREGIN07,BISTC405DCUBISTMODEREGIN08,
     BISTC405DCUBISTMODEREGIN09,BISTC405DCUBISTMODEREGIN10,BISTC405DCUBISTMODEREGIN11,
     BISTC405DCUBISTMODEREGIN12,BISTC405DCUBISTMODEREGIN13,BISTC405DCUBISTMODEREGIN14,
     BISTC405DCUBISTMODEREGIN15,BISTC405DCUBISTMODEREGIN16,BISTC405DCUBISTMODEREGIN17,
     BISTC405DCUBISTMODEREGIN18};
wire [18:0]  dcu_bist_mode_reg_out;
output     C405BISTDCUBISTMODEREGOUT00,C405BISTDCUBISTMODEREGOUT01,C405BISTDCUBISTMODEREGOUT02,
     C405BISTDCUBISTMODEREGOUT03,C405BISTDCUBISTMODEREGOUT04,C405BISTDCUBISTMODEREGOUT05,
     C405BISTDCUBISTMODEREGOUT06,C405BISTDCUBISTMODEREGOUT07,C405BISTDCUBISTMODEREGOUT08,
     C405BISTDCUBISTMODEREGOUT09,C405BISTDCUBISTMODEREGOUT10,C405BISTDCUBISTMODEREGOUT11,
     C405BISTDCUBISTMODEREGOUT12,C405BISTDCUBISTMODEREGOUT13,C405BISTDCUBISTMODEREGOUT14,
     C405BISTDCUBISTMODEREGOUT15,C405BISTDCUBISTMODEREGOUT16,C405BISTDCUBISTMODEREGOUT17,
     C405BISTDCUBISTMODEREGOUT18;
assign  {
     C405BISTDCUBISTMODEREGOUT00,C405BISTDCUBISTMODEREGOUT01,C405BISTDCUBISTMODEREGOUT02,
     C405BISTDCUBISTMODEREGOUT03,C405BISTDCUBISTMODEREGOUT04,C405BISTDCUBISTMODEREGOUT05,
     C405BISTDCUBISTMODEREGOUT06,C405BISTDCUBISTMODEREGOUT07,C405BISTDCUBISTMODEREGOUT08,
     C405BISTDCUBISTMODEREGOUT09,C405BISTDCUBISTMODEREGOUT10,C405BISTDCUBISTMODEREGOUT11,
     C405BISTDCUBISTMODEREGOUT12,C405BISTDCUBISTMODEREGOUT13,C405BISTDCUBISTMODEREGOUT14,
     C405BISTDCUBISTMODEREGOUT15,C405BISTDCUBISTMODEREGOUT16,C405BISTDCUBISTMODEREGOUT17,
     C405BISTDCUBISTMODEREGOUT18} = dcu_bist_mode_reg_out;

input          BISTC405ICUBISTMBRUN;

//input  [3:0]   BISTC405ICUBISTDEBUGSI;
wire  [3:0]   icu_bist_debug_si;
input     BISTC405ICUBISTDEBUGSI00;
input     BISTC405ICUBISTDEBUGSI01;
input     BISTC405ICUBISTDEBUGSI02;
input     BISTC405ICUBISTDEBUGSI03;
assign icu_bist_debug_si = {BISTC405ICUBISTDEBUGSI00, BISTC405ICUBISTDEBUGSI01,BISTC405ICUBISTDEBUGSI02,BISTC405ICUBISTDEBUGSI03}; 
//input  [3:0]   BISTC405ICUBISTDEBUGEN;
wire  [3:0]   icu_bist_debug_en;
input    BISTC405ICUBISTDEBUGEN00;
input    BISTC405ICUBISTDEBUGEN01;
input    BISTC405ICUBISTDEBUGEN02;
input    BISTC405ICUBISTDEBUGEN03;
assign icu_bist_debug_en = { BISTC405ICUBISTDEBUGEN00, BISTC405ICUBISTDEBUGEN01, BISTC405ICUBISTDEBUGEN02, BISTC405ICUBISTDEBUGEN03};
//output [3:0]   C405BISTICUBISTDEBUGSO;
wire [3:0]   icu_bist_debug_so;
output   C405BISTICUBISTDEBUGSO00;
output   C405BISTICUBISTDEBUGSO01;
output   C405BISTICUBISTDEBUGSO02;
output   C405BISTICUBISTDEBUGSO03;
assign {C405BISTICUBISTDEBUGSO00, C405BISTICUBISTDEBUGSO01,C405BISTICUBISTDEBUGSO02,C405BISTICUBISTDEBUGSO03} = icu_bist_debug_so ;

input          BISTC405ICUBISTSHIFTDR;
input          BISTC405ICUBISTMODEREGSI;
output         C405BISTICUBISTMODEREGSO;

input          BISTC405ICUBISTPARALLELDR;
input     BISTC405ICUBISTMODEREGIN00,BISTC405ICUBISTMODEREGIN01,BISTC405ICUBISTMODEREGIN02,
     BISTC405ICUBISTMODEREGIN03,BISTC405ICUBISTMODEREGIN04,BISTC405ICUBISTMODEREGIN05,
     BISTC405ICUBISTMODEREGIN06,BISTC405ICUBISTMODEREGIN07,BISTC405ICUBISTMODEREGIN08,
     BISTC405ICUBISTMODEREGIN09,BISTC405ICUBISTMODEREGIN10,BISTC405ICUBISTMODEREGIN11,
     BISTC405ICUBISTMODEREGIN12,BISTC405ICUBISTMODEREGIN13,BISTC405ICUBISTMODEREGIN14,
     BISTC405ICUBISTMODEREGIN15,BISTC405ICUBISTMODEREGIN16,BISTC405ICUBISTMODEREGIN17,
     BISTC405ICUBISTMODEREGIN18;
wire  [18:0]  icu_bist_mode_reg_in;
assign icu_bist_mode_reg_in = {
     BISTC405ICUBISTMODEREGIN00,BISTC405ICUBISTMODEREGIN01,BISTC405ICUBISTMODEREGIN02,
     BISTC405ICUBISTMODEREGIN03,BISTC405ICUBISTMODEREGIN04,BISTC405ICUBISTMODEREGIN05,
     BISTC405ICUBISTMODEREGIN06,BISTC405ICUBISTMODEREGIN07,BISTC405ICUBISTMODEREGIN08,
     BISTC405ICUBISTMODEREGIN09,BISTC405ICUBISTMODEREGIN10,BISTC405ICUBISTMODEREGIN11,
     BISTC405ICUBISTMODEREGIN12,BISTC405ICUBISTMODEREGIN13,BISTC405ICUBISTMODEREGIN14,
     BISTC405ICUBISTMODEREGIN15,BISTC405ICUBISTMODEREGIN16,BISTC405ICUBISTMODEREGIN17,
     BISTC405ICUBISTMODEREGIN18};
wire [18:0]  icu_bist_mode_reg_out;
output     C405BISTICUBISTMODEREGOUT00,C405BISTICUBISTMODEREGOUT01,C405BISTICUBISTMODEREGOUT02,
     C405BISTICUBISTMODEREGOUT03,C405BISTICUBISTMODEREGOUT04,C405BISTICUBISTMODEREGOUT05,
     C405BISTICUBISTMODEREGOUT06,C405BISTICUBISTMODEREGOUT07,C405BISTICUBISTMODEREGOUT08,
     C405BISTICUBISTMODEREGOUT09,C405BISTICUBISTMODEREGOUT10,C405BISTICUBISTMODEREGOUT11,
     C405BISTICUBISTMODEREGOUT12,C405BISTICUBISTMODEREGOUT13,C405BISTICUBISTMODEREGOUT14,
     C405BISTICUBISTMODEREGOUT15,C405BISTICUBISTMODEREGOUT16,C405BISTICUBISTMODEREGOUT17,
     C405BISTICUBISTMODEREGOUT18;

assign  {
     C405BISTICUBISTMODEREGOUT00,C405BISTICUBISTMODEREGOUT01,C405BISTICUBISTMODEREGOUT02,
     C405BISTICUBISTMODEREGOUT03,C405BISTICUBISTMODEREGOUT04,C405BISTICUBISTMODEREGOUT05,
     C405BISTICUBISTMODEREGOUT06,C405BISTICUBISTMODEREGOUT07,C405BISTICUBISTMODEREGOUT08,
     C405BISTICUBISTMODEREGOUT09,C405BISTICUBISTMODEREGOUT10,C405BISTICUBISTMODEREGOUT11,
     C405BISTICUBISTMODEREGOUT12,C405BISTICUBISTMODEREGOUT13,C405BISTICUBISTMODEREGOUT14,
     C405BISTICUBISTMODEREGOUT15,C405BISTICUBISTMODEREGOUT16,C405BISTICUBISTMODEREGOUT17,
     C405BISTICUBISTMODEREGOUT18} = icu_bist_mode_reg_out ;


p405s_core_top
 core(
              .C405_jtgCaptureDR(               C405JTGCAPTUREDR),
              .C405_jtgExtest(                  C405JTGEXTEST),
              .C405_jtgPgmOut(                  C405JTGPGMOUT),
              .C405_jtgShiftDR(                 C405JTGSHIFTDR),
              .C405_jtgTDO(                     C405JTGTDO),
              .C405_jtgTDOEn(                   C405JTGTDOEN),
              .C405_jtgUpdateDR(                C405JTGUPDATEDR),
              .C405_lssdDiagBistDone(           C405TESTDIAGABISTDONE),
              .C405_rstChipResetReq(            C405RSTCHIPRESETREQ),
              .C405_rstCoreResetReq(            C405RSTCORERESETREQ),
              .C405_rstSystemResetReq(          C405RSTSYSTEMRESETREQ),
              .CPU_TEType(                      {C405TRCTRIGGEREVENTTYPE0,
                                                 C405TRCTRIGGEREVENTTYPE1,
                                                 C405TRCTRIGGEREVENTTYPE2,
                                                 C405TRCTRIGGEREVENTTYPE3,
                                                 C405TRCTRIGGEREVENTTYPE4,
                                                 C405TRCTRIGGEREVENTTYPE5,
                                                 C405TRCTRIGGEREVENTTYPE6,
                                                 C405TRCTRIGGEREVENTTYPE7,
                                                 C405TRCTRIGGEREVENTTYPE8,
                                                 C405TRCTRIGGEREVENTTYPE9,
                                                 C405TRCTRIGGEREVENTTYPE10}),
              .DCS_plbABus(                     {C405PLBDCUABUS00,
                                                 C405PLBDCUABUS01,
                                                 C405PLBDCUABUS02,
                                                 C405PLBDCUABUS03,
                                                 C405PLBDCUABUS04,
                                                 C405PLBDCUABUS05,
                                                 C405PLBDCUABUS06,
                                                 C405PLBDCUABUS07,
                                                 C405PLBDCUABUS08,
                                                 C405PLBDCUABUS09,
                                                 C405PLBDCUABUS10,
                                                 C405PLBDCUABUS11,
                                                 C405PLBDCUABUS12,
                                                 C405PLBDCUABUS13,
                                                 C405PLBDCUABUS14,
                                                 C405PLBDCUABUS15,
                                                 C405PLBDCUABUS16,
                                                 C405PLBDCUABUS17,
                                                 C405PLBDCUABUS18,
                                                 C405PLBDCUABUS19,
                                                 C405PLBDCUABUS20,
                                                 C405PLBDCUABUS21,
                                                 C405PLBDCUABUS22,
                                                 C405PLBDCUABUS23,
                                                 C405PLBDCUABUS24,
                                                 C405PLBDCUABUS25,
                                                 C405PLBDCUABUS26,
                                                 C405PLBDCUABUS27,
                                                 C405PLBDCUABUS28,
                                                 C405PLBDCUABUS29,
                                                 C405PLBDCUABUS30,
                                                 C405PLBDCUABUS31}),
              .DCS_plbWrDBus(                   {C405PLBDCUWRDBUS00,
                                                 C405PLBDCUWRDBUS01,
                                                 C405PLBDCUWRDBUS02,
                                                 C405PLBDCUWRDBUS03,
                                                 C405PLBDCUWRDBUS04,
                                                 C405PLBDCUWRDBUS05,
                                                 C405PLBDCUWRDBUS06,
                                                 C405PLBDCUWRDBUS07,
                                                 C405PLBDCUWRDBUS08,
                                                 C405PLBDCUWRDBUS09,
                                                 C405PLBDCUWRDBUS10,
                                                 C405PLBDCUWRDBUS11,
                                                 C405PLBDCUWRDBUS12,
                                                 C405PLBDCUWRDBUS13,
                                                 C405PLBDCUWRDBUS14,
                                                 C405PLBDCUWRDBUS15,
                                                 C405PLBDCUWRDBUS16,
                                                 C405PLBDCUWRDBUS17,
                                                 C405PLBDCUWRDBUS18,
                                                 C405PLBDCUWRDBUS19,
                                                 C405PLBDCUWRDBUS20,
                                                 C405PLBDCUWRDBUS21,
                                                 C405PLBDCUWRDBUS22,
                                                 C405PLBDCUWRDBUS23,
                                                 C405PLBDCUWRDBUS24,
                                                 C405PLBDCUWRDBUS25,
                                                 C405PLBDCUWRDBUS26,
                                                 C405PLBDCUWRDBUS27,
                                                 C405PLBDCUWRDBUS28,
                                                 C405PLBDCUWRDBUS29,
                                                 C405PLBDCUWRDBUS30,
                                                 C405PLBDCUWRDBUS31,
                                                 C405PLBDCUWRDBUS32,
                                                 C405PLBDCUWRDBUS33,
                                                 C405PLBDCUWRDBUS34,
                                                 C405PLBDCUWRDBUS35,
                                                 C405PLBDCUWRDBUS36,
                                                 C405PLBDCUWRDBUS37,
                                                 C405PLBDCUWRDBUS38,
                                                 C405PLBDCUWRDBUS39,
                                                 C405PLBDCUWRDBUS40,
                                                 C405PLBDCUWRDBUS41,
                                                 C405PLBDCUWRDBUS42,
                                                 C405PLBDCUWRDBUS43,
                                                 C405PLBDCUWRDBUS44,
                                                 C405PLBDCUWRDBUS45,
                                                 C405PLBDCUWRDBUS46,
                                                 C405PLBDCUWRDBUS47,
                                                 C405PLBDCUWRDBUS48,
                                                 C405PLBDCUWRDBUS49,
                                                 C405PLBDCUWRDBUS50,
                                                 C405PLBDCUWRDBUS51,
                                                 C405PLBDCUWRDBUS52,
                                                 C405PLBDCUWRDBUS53,
                                                 C405PLBDCUWRDBUS54,
                                                 C405PLBDCUWRDBUS55,
                                                 C405PLBDCUWRDBUS56,
                                                 C405PLBDCUWRDBUS57,
                                                 C405PLBDCUWRDBUS58,
                                                 C405PLBDCUWRDBUS59,
                                                 C405PLBDCUWRDBUS60,
                                                 C405PLBDCUWRDBUS61,
                                                 C405PLBDCUWRDBUS62,
                                                 C405PLBDCUWRDBUS63}),
              .DCS_plbPriority(                 {C405PLBDCUPRIORITY0,
                                                 C405PLBDCUPRIORITY1}),
              .DCS_plbRNW(                      C405PLBDCURNW),
              .DCS_plbAbort(                    C405PLBDCUABORT),
              .DCU_apuWbByteEn(                 {C405APUWBBYTEEN0,
                                                 C405APUWBBYTEEN1,
                                                 C405APUWBBYTEEN2,
                                                 C405APUWBBYTEEN3}),
              .DCS_plbCacheable(                C405PLBDCUCACHEABLE),
              .DCS_plbBE(                       {C405PLBDCUBE0,
                                                 C405PLBDCUBE1,
                                                 C405PLBDCUBE2,
                                                 C405PLBDCUBE3,
                                                 C405PLBDCUBE4,
                                                 C405PLBDCUBE5,
                                                 C405PLBDCUBE6,
                                                 C405PLBDCUBE7}),
              .DCS_plbGuarded(                  C405PLBDCUGUARDED),
              .DCS_plbU0Attr(                   C405PLBDCUU0ATTR),
              .DCU_ocmAbort(                    C405DSOCMABORTOP),
              .DCU_ocmAbortReq(                 C405DSOCMABORTREQ),
              .DCU_ocmData(                     {C405DSOCMWRDBUS00,
                                                 C405DSOCMWRDBUS01,
                                                 C405DSOCMWRDBUS02,
                                                 C405DSOCMWRDBUS03,
                                                 C405DSOCMWRDBUS04,
                                                 C405DSOCMWRDBUS05,
                                                 C405DSOCMWRDBUS06,
                                                 C405DSOCMWRDBUS07,
                                                 C405DSOCMWRDBUS08,
                                                 C405DSOCMWRDBUS09,
                                                 C405DSOCMWRDBUS10,
                                                 C405DSOCMWRDBUS11,
                                                 C405DSOCMWRDBUS12,
                                                 C405DSOCMWRDBUS13,
                                                 C405DSOCMWRDBUS14,
                                                 C405DSOCMWRDBUS15,
                                                 C405DSOCMWRDBUS16,
                                                 C405DSOCMWRDBUS17,
                                                 C405DSOCMWRDBUS18,
                                                 C405DSOCMWRDBUS19,
                                                 C405DSOCMWRDBUS20,
                                                 C405DSOCMWRDBUS21,
                                                 C405DSOCMWRDBUS22,
                                                 C405DSOCMWRDBUS23,
                                                 C405DSOCMWRDBUS24,
                                                 C405DSOCMWRDBUS25,
                                                 C405DSOCMWRDBUS26,
                                                 C405DSOCMWRDBUS27,
                                                 C405DSOCMWRDBUS28,
                                                 C405DSOCMWRDBUS29,
                                                 C405DSOCMWRDBUS30,
                                                 C405DSOCMWRDBUS31}),
              .DCU_ocmLoadReq(                  C405DSOCMLOADREQ),
              .DCU_ocmStoreReq(                 C405DSOCMSTOREREQ),
              .DCU_ocmWait(                     C405DSOCMWAIT),
              .DCS_plbRequest(                  C405PLBDCUREQUEST),
              .DCS_plbSize2(                    C405PLBDCUSIZE2),
              .DCS_plbWriteThru(                C405PLBDCUWRITETHRU),
              .EXE_apuLoadData(                 {C405APUEXELOADDBUS00,
                                                 C405APUEXELOADDBUS01,
                                                 C405APUEXELOADDBUS02,
                                                 C405APUEXELOADDBUS03,
                                                 C405APUEXELOADDBUS04,
                                                 C405APUEXELOADDBUS05,
                                                 C405APUEXELOADDBUS06,
                                                 C405APUEXELOADDBUS07,
                                                 C405APUEXELOADDBUS08,
                                                 C405APUEXELOADDBUS09,
                                                 C405APUEXELOADDBUS10,
                                                 C405APUEXELOADDBUS11,
                                                 C405APUEXELOADDBUS12,
                                                 C405APUEXELOADDBUS13,
                                                 C405APUEXELOADDBUS14,
                                                 C405APUEXELOADDBUS15,
                                                 C405APUEXELOADDBUS16,
                                                 C405APUEXELOADDBUS17,
                                                 C405APUEXELOADDBUS18,
                                                 C405APUEXELOADDBUS19,
                                                 C405APUEXELOADDBUS20,
                                                 C405APUEXELOADDBUS21,
                                                 C405APUEXELOADDBUS22,
                                                 C405APUEXELOADDBUS23,
                                                 C405APUEXELOADDBUS24,
                                                 C405APUEXELOADDBUS25,
                                                 C405APUEXELOADDBUS26,
                                                 C405APUEXELOADDBUS27,
                                                 C405APUEXELOADDBUS28,
                                                 C405APUEXELOADDBUS29,
                                                 C405APUEXELOADDBUS30,
                                                 C405APUEXELOADDBUS31}),
              .EXE_dcrAddr(                     {C405DCRABUS0,
                                                 C405DCRABUS1,
                                                 C405DCRABUS2,
                                                 C405DCRABUS3,
                                                 C405DCRABUS4,
                                                 C405DCRABUS5,
                                                 C405DCRABUS6,
                                                 C405DCRABUS7,
                                                 C405DCRABUS8,
                                                 C405DCRABUS9}),
              .EXE_dcrDataBus(                  {C405DCRDBUSOUT00,
                                                 C405DCRDBUSOUT01,
                                                 C405DCRDBUSOUT02,
                                                 C405DCRDBUSOUT03,
                                                 C405DCRDBUSOUT04,
                                                 C405DCRDBUSOUT05,
                                                 C405DCRDBUSOUT06,
                                                 C405DCRDBUSOUT07,
                                                 C405DCRDBUSOUT08,
                                                 C405DCRDBUSOUT09,
                                                 C405DCRDBUSOUT10,
                                                 C405DCRDBUSOUT11,
                                                 C405DCRDBUSOUT12,
                                                 C405DCRDBUSOUT13,
                                                 C405DCRDBUSOUT14,
                                                 C405DCRDBUSOUT15,
                                                 C405DCRDBUSOUT16,
                                                 C405DCRDBUSOUT17,
                                                 C405DCRDBUSOUT18,
                                                 C405DCRDBUSOUT19,
                                                 C405DCRDBUSOUT20,
                                                 C405DCRDBUSOUT21,
                                                 C405DCRDBUSOUT22,
                                                 C405DCRDBUSOUT23,
                                                 C405DCRDBUSOUT24,
                                                 C405DCRDBUSOUT25,
                                                 C405DCRDBUSOUT26,
                                                 C405DCRDBUSOUT27,
                                                 C405DCRDBUSOUT28,
                                                 C405DCRDBUSOUT29,
                                                 C405DCRDBUSOUT30,
                                                 C405DCRDBUSOUT31}),
              .EXE_raData(                      {C405APUEXERADATA00,
                                                 C405APUEXERADATA01,
                                                 C405APUEXERADATA02,
                                                 C405APUEXERADATA03,
                                                 C405APUEXERADATA04,
                                                 C405APUEXERADATA05,
                                                 C405APUEXERADATA06,
                                                 C405APUEXERADATA07,
                                                 C405APUEXERADATA08,
                                                 C405APUEXERADATA09,
                                                 C405APUEXERADATA10,
                                                 C405APUEXERADATA11,
                                                 C405APUEXERADATA12,
                                                 C405APUEXERADATA13,
                                                 C405APUEXERADATA14,
                                                 C405APUEXERADATA15,
                                                 C405APUEXERADATA16,
                                                 C405APUEXERADATA17,
                                                 C405APUEXERADATA18,
                                                 C405APUEXERADATA19,
                                                 C405APUEXERADATA20,
                                                 C405APUEXERADATA21,
                                                 C405APUEXERADATA22,
                                                 C405APUEXERADATA23,
                                                 C405APUEXERADATA24,
                                                 C405APUEXERADATA25,
                                                 C405APUEXERADATA26,
                                                 C405APUEXERADATA27,
                                                 C405APUEXERADATA28,
                                                 C405APUEXERADATA29,
                                                 C405APUEXERADATA30,
                                                 C405APUEXERADATA31}),
              .EXE_rbData(                      {C405APUEXERBDATA00,
                                                 C405APUEXERBDATA01,
                                                 C405APUEXERBDATA02,
                                                 C405APUEXERBDATA03,
                                                 C405APUEXERBDATA04,
                                                 C405APUEXERBDATA05,
                                                 C405APUEXERBDATA06,
                                                 C405APUEXERBDATA07,
                                                 C405APUEXERBDATA08,
                                                 C405APUEXERBDATA09,
                                                 C405APUEXERBDATA10,
                                                 C405APUEXERBDATA11,
                                                 C405APUEXERBDATA12,
                                                 C405APUEXERBDATA13,
                                                 C405APUEXERBDATA14,
                                                 C405APUEXERBDATA15,
                                                 C405APUEXERBDATA16,
                                                 C405APUEXERBDATA17,
                                                 C405APUEXERBDATA18,
                                                 C405APUEXERBDATA19,
                                                 C405APUEXERBDATA20,
                                                 C405APUEXERBDATA21,
                                                 C405APUEXERBDATA22,
                                                 C405APUEXERBDATA23,
                                                 C405APUEXERBDATA24,
                                                 C405APUEXERBDATA25,
                                                 C405APUEXERBDATA26,
                                                 C405APUEXERBDATA27,
                                                 C405APUEXERBDATA28,
                                                 C405APUEXERBDATA29,
                                                 C405APUEXERBDATA30,
                                                 C405APUEXERBDATA31}),
              .EXE_xerCa(                       C405APUXERCA),
              .ICS_plbABus(                     {C405PLBICUABUS00,
                                                 C405PLBICUABUS01,
                                                 C405PLBICUABUS02,
                                                 C405PLBICUABUS03,
                                                 C405PLBICUABUS04,
                                                 C405PLBICUABUS05,
                                                 C405PLBICUABUS06,
                                                 C405PLBICUABUS07,
                                                 C405PLBICUABUS08,
                                                 C405PLBICUABUS09,
                                                 C405PLBICUABUS10,
                                                 C405PLBICUABUS11,
                                                 C405PLBICUABUS12,
                                                 C405PLBICUABUS13,
                                                 C405PLBICUABUS14,
                                                 C405PLBICUABUS15,
                                                 C405PLBICUABUS16,
                                                 C405PLBICUABUS17,
                                                 C405PLBICUABUS18,
                                                 C405PLBICUABUS19,
                                                 C405PLBICUABUS20,
                                                 C405PLBICUABUS21,
                                                 C405PLBICUABUS22,
                                                 C405PLBICUABUS23,
                                                 C405PLBICUABUS24,
                                                 C405PLBICUABUS25,
                                                 C405PLBICUABUS26,
                                                 C405PLBICUABUS27,
                                                 C405PLBICUABUS28,
                                                 C405PLBICUABUS29}),
              .ICS_plbPriority(                 {C405PLBICUPRIORITY0,
                                                 C405PLBICUPRIORITY1}),
              .ICS_plbAbort(                    C405PLBICUABORT),
              .ICS_plbCacheable(                C405PLBICUCACHEABLE),
              .ICU_ocmIcuReady(                 C405ISOCMICUREADY),
              .ICU_ocmReqPending(               C405ISOCMREQPENDING),
              .ICS_plbU0Attr(                   C405PLBICUU0ATTR),
              .ICS_plbRequest(                  C405PLBICUREQUEST),
              .ICS_plbTranSize(                 {C405PLBICUSIZE2,
                                                 C405PLBICUSIZE3}),
              .IFB_TE(                          C405TRCTRIGGEREVENTOUT),
              .IFB_cntxSyncOCM(                 C405ISOCMCONTEXTSYNC),
              .IFB_coreSleepReq(                C405CPMCORESLEEPREQ),
              .IFB_dcdFullApuL2(                C405APUDCDFULL),
              .IFB_extStopAck(                  C405DBGSTOPACK),
              .IFB_isOcmAbus(                   {C405ISOCMABUS00,
                                                 C405ISOCMABUS01,
                                                 C405ISOCMABUS02,
                                                 C405ISOCMABUS03,
                                                 C405ISOCMABUS04,
                                                 C405ISOCMABUS05,
                                                 C405ISOCMABUS06,
                                                 C405ISOCMABUS07,
                                                 C405ISOCMABUS08,
                                                 C405ISOCMABUS09,
                                                 C405ISOCMABUS10,
                                                 C405ISOCMABUS11,
                                                 C405ISOCMABUS12,
                                                 C405ISOCMABUS13,
                                                 C405ISOCMABUS14,
                                                 C405ISOCMABUS15,
                                                 C405ISOCMABUS16,
                                                 C405ISOCMABUS17,
                                                 C405ISOCMABUS18,
                                                 C405ISOCMABUS19,
                                                 C405ISOCMABUS20,
                                                 C405ISOCMABUS21,
                                                 C405ISOCMABUS22,
                                                 C405ISOCMABUS23,
                                                 C405ISOCMABUS24,
                                                 C405ISOCMABUS25,
                                                 C405ISOCMABUS26,
                                                 C405ISOCMABUS27,
                                                 C405ISOCMABUS28,
                                                 C405ISOCMABUS29}),
              .IFB_ocmAbort(                    C405ISOCMABORT),
              .IFB_reqDcdApuL2(                 {C405APUDCDINSTRUCTION00,
                                                 C405APUDCDINSTRUCTION01,
                                                 C405APUDCDINSTRUCTION02,
                                                 C405APUDCDINSTRUCTION03,
                                                 C405APUDCDINSTRUCTION04,
                                                 C405APUDCDINSTRUCTION05,
                                                 C405APUDCDINSTRUCTION06,
                                                 C405APUDCDINSTRUCTION07,
                                                 C405APUDCDINSTRUCTION08,
                                                 C405APUDCDINSTRUCTION09,
                                                 C405APUDCDINSTRUCTION10,
                                                 C405APUDCDINSTRUCTION11,
                                                 C405APUDCDINSTRUCTION12,
                                                 C405APUDCDINSTRUCTION13,
                                                 C405APUDCDINSTRUCTION14,
                                                 C405APUDCDINSTRUCTION15,
                                                 C405APUDCDINSTRUCTION16,
                                                 C405APUDCDINSTRUCTION17,
                                                 C405APUDCDINSTRUCTION18,
                                                 C405APUDCDINSTRUCTION19,
                                                 C405APUDCDINSTRUCTION20,
                                                 C405APUDCDINSTRUCTION21,
                                                 C405APUDCDINSTRUCTION22,
                                                 C405APUDCDINSTRUCTION23,
                                                 C405APUDCDINSTRUCTION24,
                                                 C405APUDCDINSTRUCTION25,
                                                 C405APUDCDINSTRUCTION26,
                                                 C405APUDCDINSTRUCTION27,
                                                 C405APUDCDINSTRUCTION28,
                                                 C405APUDCDINSTRUCTION29,
                                                 C405APUDCDINSTRUCTION30,
                                                 C405APUDCDINSTRUCTION31}),
              .IFB_wbIar(                       {C405DBGWBIAR00,
                                                 C405DBGWBIAR01,
                                                 C405DBGWBIAR02,
                                                 C405DBGWBIAR03,
                                                 C405DBGWBIAR04,
                                                 C405DBGWBIAR05,
                                                 C405DBGWBIAR06,
                                                 C405DBGWBIAR07,
                                                 C405DBGWBIAR08,
                                                 C405DBGWBIAR09,
                                                 C405DBGWBIAR10,
                                                 C405DBGWBIAR11,
                                                 C405DBGWBIAR12,
                                                 C405DBGWBIAR13,
                                                 C405DBGWBIAR14,
                                                 C405DBGWBIAR15,
                                                 C405DBGWBIAR16,
                                                 C405DBGWBIAR17,
                                                 C405DBGWBIAR18,
                                                 C405DBGWBIAR19,
                                                 C405DBGWBIAR20,
                                                 C405DBGWBIAR21,
                                                 C405DBGWBIAR22,
                                                 C405DBGWBIAR23,
                                                 C405DBGWBIAR24,
                                                 C405DBGWBIAR25,
                                                 C405DBGWBIAR26,
                                                 C405DBGWBIAR27,
                                                 C405DBGWBIAR28,
                                                 C405DBGWBIAR29}),
              .MMU_apuWbEndian(                 C405APUWBENDIAN),
              .MMU_dsocmABus(                   {C405DSOCMABUS00,
                                                 C405DSOCMABUS01,
                                                 C405DSOCMABUS02,
                                                 C405DSOCMABUS03,
                                                 C405DSOCMABUS04,
                                                 C405DSOCMABUS05,
                                                 C405DSOCMABUS06,
                                                 C405DSOCMABUS07,
                                                 C405DSOCMABUS08,
                                                 C405DSOCMABUS09,
                                                 C405DSOCMABUS10,
                                                 C405DSOCMABUS11,
                                                 C405DSOCMABUS12,
                                                 C405DSOCMABUS13,
                                                 C405DSOCMABUS14,
                                                 C405DSOCMABUS15,
                                                 C405DSOCMABUS16,
                                                 C405DSOCMABUS17,
                                                 C405DSOCMABUS18,
                                                 C405DSOCMABUS19,
                                                 C405DSOCMABUS20,
                                                 C405DSOCMABUS21,
                                                 C405DSOCMABUS22,
                                                 C405DSOCMABUS23,
                                                 C405DSOCMABUS24,
                                                 C405DSOCMABUS25,
                                                 C405DSOCMABUS26,
                                                 C405DSOCMABUS27,
                                                 C405DSOCMABUS28,
                                                 C405DSOCMABUS29}),
              .MMU_dsocmCacheable(              C405DSOCMCACHEABLE),
              .MMU_dsocmGuarded(                C405DSOCMGUARDED),
              .MMU_dsocmU0Attr(                 C405DSOCMU0ATTR),
              .MMU_dsocmXltValid(               C405DSOCMXLATEVALID),
              .MMU_isocmCacheable(              C405ISOCMCACHEABLE),
              .MMU_isocmU0Attr(                 C405ISOCMU0ATTR),
              .MMU_isocmXltValid(               C405ISOCMXLATEVALID),
              .PCL_apuExeWdCnt(                 {C405APUEXEWDCNT0,
                                                 C405APUEXEWDCNT1}),
              .PCL_apuLoadDV(                   C405APUEXELOADDVALID),
              .PCL_apuWbHold(                   C405APUWBHOLD),
              .PCL_dcdHoldForApu(               C405APUDCDHOLD),
              .PCL_dsOcmByteEn(                 {C405DSOCMBYTEEN0,
                                                 C405DSOCMBYTEEN1,
                                                 C405DSOCMBYTEEN2,
                                                 C405DSOCMBYTEEN3}),
              .PCL_exeFlushForApu(              C405APUEXEFLUSH),
              .PCL_exeHoldForApu(               C405APUEXEHOLD),
              .PCL_exeStringMultiple(           C405DSOCMSTRINGMULTIPLE),
              .PCL_mfDCR(                       C405DCRREAD),
              .PCL_mtDCR(                       C405DCRWRITE),
              .PCL_trcLoadDV(                   C405DBGLOADDATAONAPUDBUS),
              .PCL_wbComplete(                  C405DBGWBCOMPLETE),
              .PCL_wbFull(                      C405DBGWBFULL),
              .TIM_timerResetL2(                C405CPMTIMERRESETREQ),
              .TRC_evenESBusL2(                 {C405TRCEVENEXECUTIONSTATUS0,
                                                 C405TRCEVENEXECUTIONSTATUS1}),
              .TRC_oddCycle(                    C405TRCCYCLE),
              .TRC_oddESBusL2(                  {C405TRCODDEXECUTIONSTATUS0,
                                                 C405TRCODDEXECUTIONSTATUS1}),
              .TRC_tsBusL2(                     {C405TRCTRACESTATUS0,
                                                 C405TRCTRACESTATUS1,
                                                 C405TRCTRACESTATUS2,
                                                 C405TRCTRACESTATUS3}),
              .VCT_apuWbFlush(                  C405APUWBFLUSH),
              .VCT_errorOut(                    C405XXXMACHINECHECK),
              .VCT_msrCE(                       C405CPMMSRCE),
              .VCT_msrEE(                       C405CPMMSREE),
              .VCT_msrFE0(                      C405APUMSRFE0),
              .VCT_msrFE1(                      C405APUMSRFE1),
              .VCT_msrWE(                       C405DBGMSRWE),
              .VCT_timerIntrp(                  C405CPMTIMERIRQ),
              .APU_dcdApuOp(                    APUC405DCDAPUOP),
              .APU_dcdExeLdDepend(              APUC405EXELDDEPEND),
              .APU_dcdForceAlgn(                APUC405DCDFORCEALGN),
              .APU_dcdForceBESteering(          APUC405DCDFORCEBESTEERING),
              .APU_dcdFpuOp(                    APUC405DCDFPUOP),
              .APU_dcdGprWr(                    APUC405DCDGPRWRITE),
              .APU_dcdLdStByte(                 APUC405DCDLDSTBYTE),
              .APU_dcdLdStDw(                   APUC405DCDLDSTDW),
              .APU_dcdLdStHw(                   APUC405DCDLDSTHW),
              .APU_dcdLdStQw(                   APUC405DCDLDSTQW),
              .APU_dcdLdStWd(                   APUC405DCDLDSTWD),
              .APU_dcdLoad(                     APUC405DCDLOAD),
              .APU_dcdLwbLdDepend(              APUC405LWBLDDEPEND),
              .APU_dcdPrivOp(                   APUC405DCDPRIVOP),
              .APU_dcdRaEn(                     APUC405DCDRAEN),
              .APU_dcdRbEn(                     APUC405DCDRBEN),
              .APU_dcdRc(                       APUC405DCDCREN),
              .APU_dcdStore(                    APUC405DCDSTORE),
              .APU_dcdTrapBE(                   APUC405DCDTRAPBE),
              .APU_dcdTrapLE(                   APUC405DCDTRAPLE),
              .APU_dcdUpdate(                   APUC405DCDUPDATE),
              .APU_dcdValidOp(                  APUC405DCDVALIDOP),
              .APU_dcdWbLdDepend(               APUC405WBLDDEPEND),
              .APU_dcdXerCAEn(                  APUC405DCDXERCAEN),
              .APU_dcdXerOVEn(                  APUC405DCDXEROVEN),
              .APU_exception(                   APUC405EXCEPTION),
              .APU_exeBlkingMco(                APUC405EXEBLOCKINGMCO),
              .APU_exeBusy(                     APUC405EXEBUSY),
              .APU_exeCa(                       APUC405EXEXERCA),
              .APU_exeCr0(                      {APUC405EXECR0,
                                                 APUC405EXECR1,
                                                 APUC405EXECR2,
                                                 APUC405EXECR3}),
              .APU_exeCrField(                  {APUC405EXECRFIELD0,
                                                 APUC405EXECRFIELD1,
                                                 APUC405EXECRFIELD2}),
              .APU_exeNonBlkingMco(             APUC405EXENONBLOCKINGMCO),
              .APU_exeOv(                       APUC405EXEXEROV),
              .APU_exeResult(                   {APUC405EXERESULT00,
                                                 APUC405EXERESULT01,
                                                 APUC405EXERESULT02,
                                                 APUC405EXERESULT03,
                                                 APUC405EXERESULT04,
                                                 APUC405EXERESULT05,
                                                 APUC405EXERESULT06,
                                                 APUC405EXERESULT07,
                                                 APUC405EXERESULT08,
                                                 APUC405EXERESULT09,
                                                 APUC405EXERESULT10,
                                                 APUC405EXERESULT11,
                                                 APUC405EXERESULT12,
                                                 APUC405EXERESULT13,
                                                 APUC405EXERESULT14,
                                                 APUC405EXERESULT15,
                                                 APUC405EXERESULT16,
                                                 APUC405EXERESULT17,
                                                 APUC405EXERESULT18,
                                                 APUC405EXERESULT19,
                                                 APUC405EXERESULT20,
                                                 APUC405EXERESULT21,
                                                 APUC405EXERESULT22,
                                                 APUC405EXERESULT23,
                                                 APUC405EXERESULT24,
                                                 APUC405EXERESULT25,
                                                 APUC405EXERESULT26,
                                                 APUC405EXERESULT27,
                                                 APUC405EXERESULT28,
                                                 APUC405EXERESULT29,
                                                 APUC405EXERESULT30,
                                                 APUC405EXERESULT31}),
              .APU_fpuException(                APUC405FPUEXCEPTION),
              .APU_sleepReq(                    APUC405SLEEPREQ),
              .C405_timerTick(                  CPMC405TIMERTICK),
              .CB(                              CPMC405CLOCK),
              .CPM_CpuEn(                       CPMC405CPUCLKENCCLK),
              .CPM_coreClkOff(                  CPMC405CORECLKINACTIVE),
              .DBG_c405DebugHalt(               DBGC405DEBUGHALT),
              .DBG_c405ExtBusHoldAck(           DBGC405EXTBUSHOLDACK),
              .EIC_critIntrp(                   EICC405CRITINPUTIRQ),
              .EIC_extIntrp(                    EICC405EXTINPUTIRQ),
              .JTG_c405BndScanTDO(              JTGC405BNDSCANTDO),
              .JTG_c405TCK(                     JTGC405TCK),
              .JTG_c405TDI(                     JTGC405TDI),
              .JTG_c405TMS(                     JTGC405TMS),
              .JTG_c405TRST_NEG(                JTGC405TRSTNEG),
              .LSSD_bistCClk(                   TESTC405BISTCCLK),
              .LSSD_coreTestEn(                 TESTC405CNTLPOINT),
              .CPM_jtgEn(                    CPMC405JTAGCLKENCCLK),
              .LSSD_testM1(                     TESTC405TESTM1),
              .LSSD_testM3(                     TESTC405TESTM3),
              .CPM_timerEn(                  CPMC405TIMERCLKENCCLK),
              .OCM_DOF(                         DSOCMC405DISOPERANDFWD),
              .OCM_dsComplete(                  DSOCMC405COMPLETE),
              .OCM_dsData(                      {DSOCMC405RDDBUS00,
                                                 DSOCMC405RDDBUS01,
                                                 DSOCMC405RDDBUS02,
                                                 DSOCMC405RDDBUS03,
                                                 DSOCMC405RDDBUS04,
                                                 DSOCMC405RDDBUS05,
                                                 DSOCMC405RDDBUS06,
                                                 DSOCMC405RDDBUS07,
                                                 DSOCMC405RDDBUS08,
                                                 DSOCMC405RDDBUS09,
                                                 DSOCMC405RDDBUS10,
                                                 DSOCMC405RDDBUS11,
                                                 DSOCMC405RDDBUS12,
                                                 DSOCMC405RDDBUS13,
                                                 DSOCMC405RDDBUS14,
                                                 DSOCMC405RDDBUS15,
                                                 DSOCMC405RDDBUS16,
                                                 DSOCMC405RDDBUS17,
                                                 DSOCMC405RDDBUS18,
                                                 DSOCMC405RDDBUS19,
                                                 DSOCMC405RDDBUS20,
                                                 DSOCMC405RDDBUS21,
                                                 DSOCMC405RDDBUS22,
                                                 DSOCMC405RDDBUS23,
                                                 DSOCMC405RDDBUS24,
                                                 DSOCMC405RDDBUS25,
                                                 DSOCMC405RDDBUS26,
                                                 DSOCMC405RDDBUS27,
                                                 DSOCMC405RDDBUS28,
                                                 DSOCMC405RDDBUS29,
                                                 DSOCMC405RDDBUS30,
                                                 DSOCMC405RDDBUS31}),
              .OCM_dsHold(                      DSOCMC405HOLD),
              .OCM_isDATA(                      {ISOCMC405RDDBUS00,
                                                 ISOCMC405RDDBUS01,
                                                 ISOCMC405RDDBUS02,
                                                 ISOCMC405RDDBUS03,
                                                 ISOCMC405RDDBUS04,
                                                 ISOCMC405RDDBUS05,
                                                 ISOCMC405RDDBUS06,
                                                 ISOCMC405RDDBUS07,
                                                 ISOCMC405RDDBUS08,
                                                 ISOCMC405RDDBUS09,
                                                 ISOCMC405RDDBUS10,
                                                 ISOCMC405RDDBUS11,
                                                 ISOCMC405RDDBUS12,
                                                 ISOCMC405RDDBUS13,
                                                 ISOCMC405RDDBUS14,
                                                 ISOCMC405RDDBUS15,
                                                 ISOCMC405RDDBUS16,
                                                 ISOCMC405RDDBUS17,
                                                 ISOCMC405RDDBUS18,
                                                 ISOCMC405RDDBUS19,
                                                 ISOCMC405RDDBUS20,
                                                 ISOCMC405RDDBUS21,
                                                 ISOCMC405RDDBUS22,
                                                 ISOCMC405RDDBUS23,
                                                 ISOCMC405RDDBUS24,
                                                 ISOCMC405RDDBUS25,
                                                 ISOCMC405RDDBUS26,
                                                 ISOCMC405RDDBUS27,
                                                 ISOCMC405RDDBUS28,
                                                 ISOCMC405RDDBUS29,
                                                 ISOCMC405RDDBUS30,
                                                 ISOCMC405RDDBUS31,
                                                 ISOCMC405RDDBUS32,
                                                 ISOCMC405RDDBUS33,
                                                 ISOCMC405RDDBUS34,
                                                 ISOCMC405RDDBUS35,
                                                 ISOCMC405RDDBUS36,
                                                 ISOCMC405RDDBUS37,
                                                 ISOCMC405RDDBUS38,
                                                 ISOCMC405RDDBUS39,
                                                 ISOCMC405RDDBUS40,
                                                 ISOCMC405RDDBUS41,
                                                 ISOCMC405RDDBUS42,
                                                 ISOCMC405RDDBUS43,
                                                 ISOCMC405RDDBUS44,
                                                 ISOCMC405RDDBUS45,
                                                 ISOCMC405RDDBUS46,
                                                 ISOCMC405RDDBUS47,
                                                 ISOCMC405RDDBUS48,
                                                 ISOCMC405RDDBUS49,
                                                 ISOCMC405RDDBUS50,
                                                 ISOCMC405RDDBUS51,
                                                 ISOCMC405RDDBUS52,
                                                 ISOCMC405RDDBUS53,
                                                 ISOCMC405RDDBUS54,
                                                 ISOCMC405RDDBUS55,
                                                 ISOCMC405RDDBUS56,
                                                 ISOCMC405RDDBUS57,
                                                 ISOCMC405RDDBUS58,
                                                 ISOCMC405RDDBUS59,
                                                 ISOCMC405RDDBUS60,
                                                 ISOCMC405RDDBUS61,
                                                 ISOCMC405RDDBUS62,
                                                 ISOCMC405RDDBUS63}),
              .OCM_isDValid(                    {ISOCMC405RDDVALID0,
                                                 ISOCMC405RDDVALID1}),
              .OCM_isHold(                      ISOCMC405HOLD),
              .PGM_coprocPresent(               TIEC405APUPRESENT),
              .PGM_dcu_DOF(                     TIEC405DISOPERANDFWD),
              .PGM_deterministicMult(           TIEC405DETERMINISTICMULT),
              .PGM_divEn(                       TIEC405APUDIVEN),
              .PGM_mmuEn(                       TIEC405MMUEN),
              .PGM_pvrBus(                      {TIEC405PVR00,
                                                 TIEC405PVR01,
                                                 TIEC405PVR02,
                                                 TIEC405PVR03,
                                                 TIEC405PVR04,
                                                 TIEC405PVR05,
                                                 TIEC405PVR06,
                                                 TIEC405PVR07,
                                                 TIEC405PVR08,
                                                 TIEC405PVR09,
                                                 TIEC405PVR10,
                                                 TIEC405PVR11,
                                                 TIEC405PVR12,
                                                 TIEC405PVR13,
                                                 TIEC405PVR14,
                                                 TIEC405PVR15,
                                                 TIEC405PVR16,
                                                 TIEC405PVR17,
                                                 TIEC405PVR18,
                                                 TIEC405PVR19,
                                                 TIEC405PVR20,
                                                 TIEC405PVR21,
                                                 TIEC405PVR22,
                                                 TIEC405PVR23,
                                                 TIEC405PVR24,
                                                 TIEC405PVR25,
                                                 TIEC405PVR26,
                                                 TIEC405PVR27,
                                                 TIEC405PVR28,
                                                 TIEC405PVR29,
                                                 TIEC405PVR30,
                                                 TIEC405PVR31}),
              .PLB_dcuAddrAck(                  PLBC405DCUADDRACK),
              .PLB_dcuBusy(                     PLBC405DCUBUSY),
              .PLB_dcuErr(                      PLBC405DCUERR),
              .PLB_dcuRdDAck(                   PLBC405DCURDDACK),
              .PLB_dcuRdDBus(                   {PLBC405DCURDDBUS00,
                                                 PLBC405DCURDDBUS01,
                                                 PLBC405DCURDDBUS02,
                                                 PLBC405DCURDDBUS03,
                                                 PLBC405DCURDDBUS04,
                                                 PLBC405DCURDDBUS05,
                                                 PLBC405DCURDDBUS06,
                                                 PLBC405DCURDDBUS07,
                                                 PLBC405DCURDDBUS08,
                                                 PLBC405DCURDDBUS09,
                                                 PLBC405DCURDDBUS10,
                                                 PLBC405DCURDDBUS11,
                                                 PLBC405DCURDDBUS12,
                                                 PLBC405DCURDDBUS13,
                                                 PLBC405DCURDDBUS14,
                                                 PLBC405DCURDDBUS15,
                                                 PLBC405DCURDDBUS16,
                                                 PLBC405DCURDDBUS17,
                                                 PLBC405DCURDDBUS18,
                                                 PLBC405DCURDDBUS19,
                                                 PLBC405DCURDDBUS20,
                                                 PLBC405DCURDDBUS21,
                                                 PLBC405DCURDDBUS22,
                                                 PLBC405DCURDDBUS23,
                                                 PLBC405DCURDDBUS24,
                                                 PLBC405DCURDDBUS25,
                                                 PLBC405DCURDDBUS26,
                                                 PLBC405DCURDDBUS27,
                                                 PLBC405DCURDDBUS28,
                                                 PLBC405DCURDDBUS29,
                                                 PLBC405DCURDDBUS30,
                                                 PLBC405DCURDDBUS31,
                                                 PLBC405DCURDDBUS32,
                                                 PLBC405DCURDDBUS33,
                                                 PLBC405DCURDDBUS34,
                                                 PLBC405DCURDDBUS35,
                                                 PLBC405DCURDDBUS36,
                                                 PLBC405DCURDDBUS37,
                                                 PLBC405DCURDDBUS38,
                                                 PLBC405DCURDDBUS39,
                                                 PLBC405DCURDDBUS40,
                                                 PLBC405DCURDDBUS41,
                                                 PLBC405DCURDDBUS42,
                                                 PLBC405DCURDDBUS43,
                                                 PLBC405DCURDDBUS44,
                                                 PLBC405DCURDDBUS45,
                                                 PLBC405DCURDDBUS46,
                                                 PLBC405DCURDDBUS47,
                                                 PLBC405DCURDDBUS48,
                                                 PLBC405DCURDDBUS49,
                                                 PLBC405DCURDDBUS50,
                                                 PLBC405DCURDDBUS51,
                                                 PLBC405DCURDDBUS52,
                                                 PLBC405DCURDDBUS53,
                                                 PLBC405DCURDDBUS54,
                                                 PLBC405DCURDDBUS55,
                                                 PLBC405DCURDDBUS56,
                                                 PLBC405DCURDDBUS57,
                                                 PLBC405DCURDDBUS58,
                                                 PLBC405DCURDDBUS59,
                                                 PLBC405DCURDDBUS60,
                                                 PLBC405DCURDDBUS61,
                                                 PLBC405DCURDDBUS62,
                                                 PLBC405DCURDDBUS63}),
              .PLB_dcuRdWdAddr(                 {PLBC405DCURDWDADDR1,
                                                 PLBC405DCURDWDADDR2,
                                                 PLBC405DCURDWDADDR3}),
              .PLB_dcuSsize(                    PLBC405DCUSSIZE1),
              .PLB_dcuWrDAck(                   PLBC405DCUWRDACK),
              .PLB_icuAddrAck(                  PLBC405ICUADDRACK),
              .PLB_icuBusy(                     PLBC405ICUBUSY),
              .PLB_icuDBus(                     {PLBC405ICURDDBUS00,
                                                 PLBC405ICURDDBUS01,
                                                 PLBC405ICURDDBUS02,
                                                 PLBC405ICURDDBUS03,
                                                 PLBC405ICURDDBUS04,
                                                 PLBC405ICURDDBUS05,
                                                 PLBC405ICURDDBUS06,
                                                 PLBC405ICURDDBUS07,
                                                 PLBC405ICURDDBUS08,
                                                 PLBC405ICURDDBUS09,
                                                 PLBC405ICURDDBUS10,
                                                 PLBC405ICURDDBUS11,
                                                 PLBC405ICURDDBUS12,
                                                 PLBC405ICURDDBUS13,
                                                 PLBC405ICURDDBUS14,
                                                 PLBC405ICURDDBUS15,
                                                 PLBC405ICURDDBUS16,
                                                 PLBC405ICURDDBUS17,
                                                 PLBC405ICURDDBUS18,
                                                 PLBC405ICURDDBUS19,
                                                 PLBC405ICURDDBUS20,
                                                 PLBC405ICURDDBUS21,
                                                 PLBC405ICURDDBUS22,
                                                 PLBC405ICURDDBUS23,
                                                 PLBC405ICURDDBUS24,
                                                 PLBC405ICURDDBUS25,
                                                 PLBC405ICURDDBUS26,
                                                 PLBC405ICURDDBUS27,
                                                 PLBC405ICURDDBUS28,
                                                 PLBC405ICURDDBUS29,
                                                 PLBC405ICURDDBUS30,
                                                 PLBC405ICURDDBUS31,
                                                 PLBC405ICURDDBUS32,
                                                 PLBC405ICURDDBUS33,
                                                 PLBC405ICURDDBUS34,
                                                 PLBC405ICURDDBUS35,
                                                 PLBC405ICURDDBUS36,
                                                 PLBC405ICURDDBUS37,
                                                 PLBC405ICURDDBUS38,
                                                 PLBC405ICURDDBUS39,
                                                 PLBC405ICURDDBUS40,
                                                 PLBC405ICURDDBUS41,
                                                 PLBC405ICURDDBUS42,
                                                 PLBC405ICURDDBUS43,
                                                 PLBC405ICURDDBUS44,
                                                 PLBC405ICURDDBUS45,
                                                 PLBC405ICURDDBUS46,
                                                 PLBC405ICURDDBUS47,
                                                 PLBC405ICURDDBUS48,
                                                 PLBC405ICURDDBUS49,
                                                 PLBC405ICURDDBUS50,
                                                 PLBC405ICURDDBUS51,
                                                 PLBC405ICURDDBUS52,
                                                 PLBC405ICURDDBUS53,
                                                 PLBC405ICURDDBUS54,
                                                 PLBC405ICURDDBUS55,
                                                 PLBC405ICURDDBUS56,
                                                 PLBC405ICURDDBUS57,
                                                 PLBC405ICURDDBUS58,
                                                 PLBC405ICURDDBUS59,
                                                 PLBC405ICURDDBUS60,
                                                 PLBC405ICURDDBUS61,
                                                 PLBC405ICURDDBUS62,
                                                 PLBC405ICURDDBUS63}),
              .PLB_icuError(                    PLBC405ICUERR),
              .PLB_icuRdDAck(                   PLBC405ICURDDACK),
              .PLB_icuRdWrAddr(                 {PLBC405ICURDWDADDR1,
                                                 PLBC405ICURDWDADDR2,
                                                 PLBC405ICURDWDADDR3}),
              .PLB_icuSSize(                    PLBC405ICUSSIZE1),
              .PLB_sampleCycle(                 CPMC405PLBSAMPLECYCLE),
              .RST_c405ResetChip(               RSTC405RESETCHIP),
              .RST_c405ResetSystem(             RSTC405RESETSYSTEM),
              .TRC_c405TE(                      TRCC405TRIGGEREVENTIN),
              .TRC_c405TraceDisable(            TRCC405TRACEDISABLE),
              .XXX_dcrAck(                      DCRC405ACK),
              .XXX_dcrDataBus(                  {DCRC405DBUSIN00,
                                                 DCRC405DBUSIN01,
                                                 DCRC405DBUSIN02,
                                                 DCRC405DBUSIN03,
                                                 DCRC405DBUSIN04,
                                                 DCRC405DBUSIN05,
                                                 DCRC405DBUSIN06,
                                                 DCRC405DBUSIN07,
                                                 DCRC405DBUSIN08,
                                                 DCRC405DBUSIN09,
                                                 DCRC405DBUSIN10,
                                                 DCRC405DBUSIN11,
                                                 DCRC405DBUSIN12,
                                                 DCRC405DBUSIN13,
                                                 DCRC405DBUSIN14,
                                                 DCRC405DBUSIN15,
                                                 DCRC405DBUSIN16,
                                                 DCRC405DBUSIN17,
                                                 DCRC405DBUSIN18,
                                                 DCRC405DBUSIN19,
                                                 DCRC405DBUSIN20,
                                                 DCRC405DBUSIN21,
                                                 DCRC405DBUSIN22,
                                                 DCRC405DBUSIN23,
                                                 DCRC405DBUSIN24,
                                                 DCRC405DBUSIN25,
                                                 DCRC405DBUSIN26,
                                                 DCRC405DBUSIN27,
                                                 DCRC405DBUSIN28,
                                                 DCRC405DBUSIN29,
                                                 DCRC405DBUSIN30,
                                                 DCRC405DBUSIN31}),
              .XXX_uncondEvent(                 DBGC405UNCONDDEBUGEVENT),
              .resetCore(                       RSTC405RESETCORE),
              .BIST_pepsPF(                     {C405BISTPEPSPF00,
                                                 C405BISTPEPSPF01,
                                                 C405BISTPEPSPF02}),
              .LSSD_c405CE0EVS(                 TESTC405CE0EVS),
              .LSSD_c405BistCE0StClk(           TESTC405BISTCE0STCLK),
              .LSSD_c405BistCE1Enable(          TESTC405BISTCE1ENABLE),
              .LSSD_c405BistCE1Mode(            TESTC405BISTCE1MODE),
              .TIE_c405ClockEnable(             TIEC405CLOCKENABLE),
              .TIE_c405DutyEnable(              TIEC405DUTYENABLE),
              .CPM_c405PLBClock(                CPMC405PLBSYNCCLOCK),
              .CPM_c405SyncBypass(              CPMC405SYNCBYPASS),
              .PLB_sampleCycleAlt(              CPMC405PLBSAMPLECYCLEALT),
              .testmode(                        TESTC405TESTMODE),
              .dcu_bist_debug_si(               dcu_bist_debug_si),  // BIST ports
              .dcu_bist_debug_so(               dcu_bist_debug_so),
              .dcu_bist_debug_en(               dcu_bist_debug_en),
              .dcu_bist_mode_reg_in(            dcu_bist_mode_reg_in),
              .dcu_bist_mode_reg_out(           dcu_bist_mode_reg_out),
              .dcu_bist_parallel_dr(            BISTC405DCUBISTPARALLELDR),
              .dcu_bist_mode_reg_si(            BISTC405DCUBISTMODEREGSI),
              .dcu_bist_mode_reg_so(            C405BISTDCUBISTMODEREGSO),
              .dcu_bist_shift_dr(               BISTC405DCUBISTSHIFTDR),
              .dcu_bist_mbrun(                  BISTC405DCUBISTMBRUN),
              .icu_bist_debug_si(               icu_bist_debug_si),
              .icu_bist_debug_so(               icu_bist_debug_so),
              .icu_bist_debug_en(               icu_bist_debug_en),
              .icu_bist_mode_reg_in(            icu_bist_mode_reg_in),
              .icu_bist_mode_reg_out(           icu_bist_mode_reg_out),
              .icu_bist_parallel_dr(            BISTC405ICUBISTPARALLELDR),
              .icu_bist_mode_reg_si(            BISTC405ICUBISTMODEREGSI),
              .icu_bist_mode_reg_so(            C405BISTICUBISTMODEREGSO),
              .icu_bist_shift_dr(               BISTC405ICUBISTSHIFTDR),
              .icu_bist_mbrun(                  BISTC405ICUBISTMBRUN)
             );

endmodule
