library verilog;
use verilog.vl_types.all;
entity t_altivec_env_pkg is
end t_altivec_env_pkg;
