library verilog;
use verilog.vl_types.all;
entity p405s_dcu_top is
    port(
        CAR_mmuAttr_E1  : out    vl_logic;
        CAR_mmuAttr_E2  : out    vl_logic;
        DCU_CA          : out    vl_logic;
        DCU_DA          : out    vl_logic;
        DCU_SCL2        : out    vl_logic;
        DCU_SDQ_mod_NEG : out    vl_logic_vector(0 to 31);
        DCU_apuWbByteEn : out    vl_logic_vector(0 to 3);
        DCU_carByteEn   : out    vl_logic_vector(0 to 3);
        DCU_data_NEG    : out    vl_logic_vector(0 to 31);
        DCU_diagBus     : out    vl_logic_vector(0 to 20);
        DCU_firstCycCarStXltV: out    vl_logic;
        DCU_icuSize     : out    vl_logic_vector(0 to 2);
        DCU_ocmAbort    : out    vl_logic;
        DCU_ocmData     : out    vl_logic_vector(0 to 31);
        DCU_ocmLoadReq  : out    vl_logic;
        DCU_ocmStoreReq : out    vl_logic;
        DCU_ocmWait     : out    vl_logic;
        DCU_pclOcmLdPendNoWait: out    vl_logic;
        DCU_plbABus     : out    vl_logic_vector(0 to 31);
        DCU_plbAbort    : out    vl_logic;
        DCU_plbCacheable: out    vl_logic;
        DCU_plbDBus     : out    vl_logic_vector(0 to 63);
        DCU_plbDTags    : out    vl_logic_vector(0 to 7);
        DCU_plbGuarded  : out    vl_logic;
        DCU_plbPriority : out    vl_logic;
        DCU_plbRNW      : out    vl_logic;
        DCU_plbRequest  : out    vl_logic;
        DCU_plbTranSize : out    vl_logic;
        DCU_plbU0Attr   : out    vl_logic;
        DCU_plbWriteThru: out    vl_logic;
        DCU_sleepReq    : out    vl_logic;
        CAR_U0Attr      : in     vl_logic;
        CAR_cacheable   : in     vl_logic;
        CAR_endian      : in     vl_logic;
        CAR_guarded     : in     vl_logic;
        CAR_writethru   : in     vl_logic;
        CB              : in     vl_logic;
        EXE_dcuData     : in     vl_logic_vector(0 to 31);
        ICU_dcuCCR0_L2  : in     vl_logic_vector(0 to 11);
        ICU_syncAfterReset: in     vl_logic;
        MMU_dcuShadowAbort: in     vl_logic;
        MMU_dcuUTLBAbort: in     vl_logic;
        MMU_dcuXltValid : in     vl_logic;
        MMU_diagOut     : in     vl_logic_vector(0 to 2);
        MMU_dsRA        : in     vl_logic_vector(0 to 29);
        MMU_wbHold      : in     vl_logic;
        OCM_dsComplete  : in     vl_logic;
        OCM_dsHold      : in     vl_logic;
        PCL_dcuByteEn   : in     vl_logic_vector(0 to 3);
        PCL_dcuOp       : in     vl_logic_vector(0 to 11);
        PCL_dcuOp_early : in     vl_logic_vector(0 to 2);
        PCL_stSteerCntl : in     vl_logic_vector(0 to 9);
        PLB_dcuAddrAck  : in     vl_logic;
        PLB_dcuBusy     : in     vl_logic;
        PLB_dcuRdDAck   : in     vl_logic;
        PLB_dcuRdDBus   : in     vl_logic_vector(0 to 63);
        PLB_dcuRdWdAddr : in     vl_logic_vector(0 to 2);
        PLB_dcuSsize    : in     vl_logic;
        PLB_dcuWrDAck   : in     vl_logic;
        PLB_sampleCycle : in     vl_logic;
        VCT_exeAbort    : in     vl_logic;
        VCT_wbAbort     : in     vl_logic;
        resetCore       : in     vl_logic;
        testEn          : in     vl_logic;
        DCU_parityError : out    vl_logic;
        DCU_FlushParityError: out    vl_logic;
        ICU_CCR1DCTE    : in     vl_logic;
        ICU_CCR1DCDE    : in     vl_logic;
        PLB_sampleCycleAlt: in     vl_logic;
        CPM_c405SyncBypass: in     vl_logic;
        dcu_bist_debug_si: in     vl_logic_vector(3 downto 0);
        dcu_bist_debug_so: out    vl_logic_vector(3 downto 0);
        dcu_bist_debug_en: in     vl_logic_vector(3 downto 0);
        dcu_bist_mode_reg_in: in     vl_logic_vector(18 downto 0);
        dcu_bist_mode_reg_out: out    vl_logic_vector(18 downto 0);
        dcu_bist_parallel_dr: in     vl_logic;
        dcu_bist_mode_reg_si: in     vl_logic;
        dcu_bist_mode_reg_so: out    vl_logic;
        dcu_bist_shift_dr: in     vl_logic;
        dcu_bist_mbrun  : in     vl_logic;
        resetMemBist    : in     vl_logic
    );
end p405s_dcu_top;
