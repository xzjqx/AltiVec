library verilog;
use verilog.vl_types.all;
entity p405s_wbStage is
    port(
        PCL_ldAdjE2     : out    vl_logic_vector(1 to 3);
        PCL_ldFillByPassMuxSel: out    vl_logic_vector(0 to 5);
        ldAdjSel        : out    vl_logic_vector(1 to 3);
        PCL_ldSteerMuxSel: out    vl_logic_vector(0 to 7);
        PCL_wbRpWrEn    : out    vl_logic;
        wbFull          : out    vl_logic;
        wbLoad          : out    vl_logic;
        wbLpWrEn        : out    vl_logic;
        CB              : in     vl_logic;
        byteCount       : in     vl_logic_vector(6 to 7);
        cntGtEq4        : in     vl_logic;
        exeAlg          : in     vl_logic;
        exeByteRev      : in     vl_logic;
        exeStorageOp    : in     vl_logic;
        exeEA           : in     vl_logic_vector(30 to 31);
        exeLoadQ        : in     vl_logic;
        exeMultiple     : in     vl_logic;
        exeRpWrEnQ      : in     vl_logic;
        exeStrgSt       : in     vl_logic_vector(0 to 2);
        exeString       : in     vl_logic;
        loadSteerMuxSel : in     vl_logic;
        lwbE1           : in     vl_logic;
        nxtWbLpWrEn     : in     vl_logic;
        PCL_wbStorageOp : out    vl_logic;
        wbClearOrFlush  : in     vl_logic;
        wbEndian        : in     vl_logic;
        wbE1            : in     vl_logic;
        wbE2            : in     vl_logic;
        wbStrgLS        : out    vl_logic;
        exeLwarx        : in     vl_logic;
        exeStwcx        : in     vl_logic;
        wbLwarx         : out    vl_logic;
        wbStwcx         : out    vl_logic;
        exeApuFpuLoad   : in     vl_logic;
        wbApuFpuLoad    : out    vl_logic;
        algnErr         : in     vl_logic;
        PCL_wbAlgnErr   : out    vl_logic;
        exeLdNotSt      : in     vl_logic;
        PCL_wbLdNotSt   : out    vl_logic;
        exeStore        : in     vl_logic;
        exeWUD          : in     vl_logic;
        wbLdOrStWUD     : out    vl_logic;
        wbStrgC1        : out    vl_logic;
        exeRA           : in     vl_logic_vector(0 to 4);
        wbRAL2          : out    vl_logic_vector(0 to 4);
        exeStrgEnd      : in     vl_logic;
        PCL_wbStrgEnd   : out    vl_logic;
        exeByteEn       : in     vl_logic_vector(0 to 3);
        wbByteEn        : out    vl_logic_vector(0 to 3);
        wbFullForPO     : out    vl_logic;
        exeTrapLE       : in     vl_logic;
        exeTrapBE       : in     vl_logic;
        exeApuFpuLdSt   : in     vl_logic;
        wbStrgSt        : out    vl_logic_vector(1 to 2);
        wbFullForDepend : out    vl_logic;
        wbLoadForApu    : out    vl_logic
    );
end p405s_wbStage;
