library verilog;
use verilog.vl_types.all;
entity p405s_sync_top is
    port(
        ICS_plbABus     : out    vl_logic_vector(0 to 29);
        ICS_plbAbort    : out    vl_logic;
        ICS_plbCacheable: out    vl_logic;
        ICS_plbRequest  : out    vl_logic;
        ICS_plbTranSize : out    vl_logic_vector(2 to 3);
        ICS_plbU0Attr   : out    vl_logic;
        ICS_plbPriority : out    vl_logic_vector(0 to 1);
        ICS_c405AddrAck : out    vl_logic;
        ICS_c405IcuBusy : out    vl_logic;
        ICS_c405Error   : out    vl_logic;
        ICS_c405RdDAck  : out    vl_logic;
        ICS_c405DBus    : out    vl_logic_vector(0 to 63);
        ICS_c405RdWrAddr: out    vl_logic_vector(1 to 3);
        ICS_c405SSize   : out    vl_logic;
        C405_icsABus    : in     vl_logic_vector(0 to 29);
        C405_icsAbort   : in     vl_logic;
        C405_icsCacheable: in     vl_logic;
        C405_icsRequest : in     vl_logic;
        C405_icsTranSize: in     vl_logic_vector(2 to 3);
        C405_icsU0Attr  : in     vl_logic;
        C405_icsPriority: in     vl_logic_vector(0 to 1);
        PLB_icsAddrAck  : in     vl_logic;
        PLB_icsIcuBusy  : in     vl_logic;
        PLB_icsError    : in     vl_logic;
        PLB_icsRdDAck   : in     vl_logic;
        PLB_icsDBus     : in     vl_logic_vector(0 to 63);
        PLB_icsRdWrAddr : in     vl_logic_vector(1 to 3);
        PLB_icsSSize    : in     vl_logic;
        DCS_plbRequest  : out    vl_logic;
        DCS_plbRNW      : out    vl_logic;
        DCS_plbABus     : out    vl_logic_vector(0 to 31);
        DCS_plbSize2    : out    vl_logic;
        DCS_plbCacheable: out    vl_logic;
        DCS_plbWriteThru: out    vl_logic;
        DCS_plbU0Attr   : out    vl_logic;
        DCS_plbGuarded  : out    vl_logic;
        DCS_plbBE       : out    vl_logic_vector(0 to 7);
        DCS_plbPriority : out    vl_logic_vector(0 to 1);
        DCS_plbAbort    : out    vl_logic;
        DCS_plbWrDBus   : out    vl_logic_vector(0 to 63);
        DCS_c405AddrAck : out    vl_logic;
        DCS_c405SSize1  : out    vl_logic;
        DCS_c405RdDAck  : out    vl_logic;
        DCS_c405RdDBus  : out    vl_logic_vector(0 to 63);
        DCS_c405RdWdAddr: out    vl_logic_vector(1 to 3);
        DCS_c405WrDAck  : out    vl_logic;
        DCS_c405Busy    : out    vl_logic;
        DCS_c405Err     : out    vl_logic;
        C405_dcsDcuRequest: in     vl_logic;
        C405_dcsDcuRNW  : in     vl_logic;
        C405_dcsDcuABus : in     vl_logic_vector(0 to 31);
        C405_dcsDcuSize2: in     vl_logic;
        C405_dcsDcuCacheable: in     vl_logic;
        C405_dcsDcuWriteThru: in     vl_logic;
        C405_dcsDcuU0Attr: in     vl_logic;
        C405_dcsDcuGuarded: in     vl_logic;
        C405_dcsDcuBE   : in     vl_logic_vector(0 to 7);
        C405_dcsDcuPriority: in     vl_logic_vector(0 to 1);
        C405_dcsDcuAbort: in     vl_logic;
        C405_dcsDcuWrDBus: in     vl_logic_vector(0 to 63);
        PLB_dcsAddrAck  : in     vl_logic;
        PLB_dcsSSize1   : in     vl_logic;
        PLB_dcsRdDAck   : in     vl_logic;
        PLB_dcsRdDBus   : in     vl_logic_vector(0 to 63);
        PLB_dcsRdWdAddr : in     vl_logic_vector(1 to 3);
        PLB_dcsWrDAck   : in     vl_logic;
        PLB_dcsBusy     : in     vl_logic;
        PLB_dcsErr      : in     vl_logic;
        CPM_c405SyncBypass: in     vl_logic;
        EXT_sysclkPLB   : in     vl_logic;
        CB              : in     vl_logic;
        RST_ResetCore   : in     vl_logic
    );
end p405s_sync_top;
