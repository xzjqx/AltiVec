library verilog;
use verilog.vl_types.all;
entity PPC405F5V1 is
    port(
        C405APUDCDFULL  : out    vl_logic;
        C405APUDCDHOLD  : out    vl_logic;
        C405APUDCDINSTRUCTION00: out    vl_logic;
        C405APUDCDINSTRUCTION01: out    vl_logic;
        C405APUDCDINSTRUCTION02: out    vl_logic;
        C405APUDCDINSTRUCTION03: out    vl_logic;
        C405APUDCDINSTRUCTION04: out    vl_logic;
        C405APUDCDINSTRUCTION05: out    vl_logic;
        C405APUDCDINSTRUCTION06: out    vl_logic;
        C405APUDCDINSTRUCTION07: out    vl_logic;
        C405APUDCDINSTRUCTION08: out    vl_logic;
        C405APUDCDINSTRUCTION09: out    vl_logic;
        C405APUDCDINSTRUCTION10: out    vl_logic;
        C405APUDCDINSTRUCTION11: out    vl_logic;
        C405APUDCDINSTRUCTION12: out    vl_logic;
        C405APUDCDINSTRUCTION13: out    vl_logic;
        C405APUDCDINSTRUCTION14: out    vl_logic;
        C405APUDCDINSTRUCTION15: out    vl_logic;
        C405APUDCDINSTRUCTION16: out    vl_logic;
        C405APUDCDINSTRUCTION17: out    vl_logic;
        C405APUDCDINSTRUCTION18: out    vl_logic;
        C405APUDCDINSTRUCTION19: out    vl_logic;
        C405APUDCDINSTRUCTION20: out    vl_logic;
        C405APUDCDINSTRUCTION21: out    vl_logic;
        C405APUDCDINSTRUCTION22: out    vl_logic;
        C405APUDCDINSTRUCTION23: out    vl_logic;
        C405APUDCDINSTRUCTION24: out    vl_logic;
        C405APUDCDINSTRUCTION25: out    vl_logic;
        C405APUDCDINSTRUCTION26: out    vl_logic;
        C405APUDCDINSTRUCTION27: out    vl_logic;
        C405APUDCDINSTRUCTION28: out    vl_logic;
        C405APUDCDINSTRUCTION29: out    vl_logic;
        C405APUDCDINSTRUCTION30: out    vl_logic;
        C405APUDCDINSTRUCTION31: out    vl_logic;
        C405APUEXEFLUSH : out    vl_logic;
        C405APUEXEHOLD  : out    vl_logic;
        C405APUEXELOADDBUS00: out    vl_logic;
        C405APUEXELOADDBUS01: out    vl_logic;
        C405APUEXELOADDBUS02: out    vl_logic;
        C405APUEXELOADDBUS03: out    vl_logic;
        C405APUEXELOADDBUS04: out    vl_logic;
        C405APUEXELOADDBUS05: out    vl_logic;
        C405APUEXELOADDBUS06: out    vl_logic;
        C405APUEXELOADDBUS07: out    vl_logic;
        C405APUEXELOADDBUS08: out    vl_logic;
        C405APUEXELOADDBUS09: out    vl_logic;
        C405APUEXELOADDBUS10: out    vl_logic;
        C405APUEXELOADDBUS11: out    vl_logic;
        C405APUEXELOADDBUS12: out    vl_logic;
        C405APUEXELOADDBUS13: out    vl_logic;
        C405APUEXELOADDBUS14: out    vl_logic;
        C405APUEXELOADDBUS15: out    vl_logic;
        C405APUEXELOADDBUS16: out    vl_logic;
        C405APUEXELOADDBUS17: out    vl_logic;
        C405APUEXELOADDBUS18: out    vl_logic;
        C405APUEXELOADDBUS19: out    vl_logic;
        C405APUEXELOADDBUS20: out    vl_logic;
        C405APUEXELOADDBUS21: out    vl_logic;
        C405APUEXELOADDBUS22: out    vl_logic;
        C405APUEXELOADDBUS23: out    vl_logic;
        C405APUEXELOADDBUS24: out    vl_logic;
        C405APUEXELOADDBUS25: out    vl_logic;
        C405APUEXELOADDBUS26: out    vl_logic;
        C405APUEXELOADDBUS27: out    vl_logic;
        C405APUEXELOADDBUS28: out    vl_logic;
        C405APUEXELOADDBUS29: out    vl_logic;
        C405APUEXELOADDBUS30: out    vl_logic;
        C405APUEXELOADDBUS31: out    vl_logic;
        C405APUEXELOADDVALID: out    vl_logic;
        C405APUEXERADATA00: out    vl_logic;
        C405APUEXERADATA01: out    vl_logic;
        C405APUEXERADATA02: out    vl_logic;
        C405APUEXERADATA03: out    vl_logic;
        C405APUEXERADATA04: out    vl_logic;
        C405APUEXERADATA05: out    vl_logic;
        C405APUEXERADATA06: out    vl_logic;
        C405APUEXERADATA07: out    vl_logic;
        C405APUEXERADATA08: out    vl_logic;
        C405APUEXERADATA09: out    vl_logic;
        C405APUEXERADATA10: out    vl_logic;
        C405APUEXERADATA11: out    vl_logic;
        C405APUEXERADATA12: out    vl_logic;
        C405APUEXERADATA13: out    vl_logic;
        C405APUEXERADATA14: out    vl_logic;
        C405APUEXERADATA15: out    vl_logic;
        C405APUEXERADATA16: out    vl_logic;
        C405APUEXERADATA17: out    vl_logic;
        C405APUEXERADATA18: out    vl_logic;
        C405APUEXERADATA19: out    vl_logic;
        C405APUEXERADATA20: out    vl_logic;
        C405APUEXERADATA21: out    vl_logic;
        C405APUEXERADATA22: out    vl_logic;
        C405APUEXERADATA23: out    vl_logic;
        C405APUEXERADATA24: out    vl_logic;
        C405APUEXERADATA25: out    vl_logic;
        C405APUEXERADATA26: out    vl_logic;
        C405APUEXERADATA27: out    vl_logic;
        C405APUEXERADATA28: out    vl_logic;
        C405APUEXERADATA29: out    vl_logic;
        C405APUEXERADATA30: out    vl_logic;
        C405APUEXERADATA31: out    vl_logic;
        C405APUEXERBDATA00: out    vl_logic;
        C405APUEXERBDATA01: out    vl_logic;
        C405APUEXERBDATA02: out    vl_logic;
        C405APUEXERBDATA03: out    vl_logic;
        C405APUEXERBDATA04: out    vl_logic;
        C405APUEXERBDATA05: out    vl_logic;
        C405APUEXERBDATA06: out    vl_logic;
        C405APUEXERBDATA07: out    vl_logic;
        C405APUEXERBDATA08: out    vl_logic;
        C405APUEXERBDATA09: out    vl_logic;
        C405APUEXERBDATA10: out    vl_logic;
        C405APUEXERBDATA11: out    vl_logic;
        C405APUEXERBDATA12: out    vl_logic;
        C405APUEXERBDATA13: out    vl_logic;
        C405APUEXERBDATA14: out    vl_logic;
        C405APUEXERBDATA15: out    vl_logic;
        C405APUEXERBDATA16: out    vl_logic;
        C405APUEXERBDATA17: out    vl_logic;
        C405APUEXERBDATA18: out    vl_logic;
        C405APUEXERBDATA19: out    vl_logic;
        C405APUEXERBDATA20: out    vl_logic;
        C405APUEXERBDATA21: out    vl_logic;
        C405APUEXERBDATA22: out    vl_logic;
        C405APUEXERBDATA23: out    vl_logic;
        C405APUEXERBDATA24: out    vl_logic;
        C405APUEXERBDATA25: out    vl_logic;
        C405APUEXERBDATA26: out    vl_logic;
        C405APUEXERBDATA27: out    vl_logic;
        C405APUEXERBDATA28: out    vl_logic;
        C405APUEXERBDATA29: out    vl_logic;
        C405APUEXERBDATA30: out    vl_logic;
        C405APUEXERBDATA31: out    vl_logic;
        C405APUEXEWDCNT0: out    vl_logic;
        C405APUEXEWDCNT1: out    vl_logic;
        C405APUMSRFE0   : out    vl_logic;
        C405APUMSRFE1   : out    vl_logic;
        C405APUWBBYTEEN0: out    vl_logic;
        C405APUWBBYTEEN1: out    vl_logic;
        C405APUWBBYTEEN2: out    vl_logic;
        C405APUWBBYTEEN3: out    vl_logic;
        C405APUWBENDIAN : out    vl_logic;
        C405APUWBFLUSH  : out    vl_logic;
        C405APUWBHOLD   : out    vl_logic;
        C405APUXERCA    : out    vl_logic;
        C405CPMCORESLEEPREQ: out    vl_logic;
        C405CPMMSRCE    : out    vl_logic;
        C405CPMMSREE    : out    vl_logic;
        C405CPMTIMERIRQ : out    vl_logic;
        C405CPMTIMERRESETREQ: out    vl_logic;
        C405DBGLOADDATAONAPUDBUS: out    vl_logic;
        C405DBGMSRWE    : out    vl_logic;
        C405DBGSTOPACK  : out    vl_logic;
        C405DBGWBCOMPLETE: out    vl_logic;
        C405DBGWBFULL   : out    vl_logic;
        C405DBGWBIAR00  : out    vl_logic;
        C405DBGWBIAR01  : out    vl_logic;
        C405DBGWBIAR02  : out    vl_logic;
        C405DBGWBIAR03  : out    vl_logic;
        C405DBGWBIAR04  : out    vl_logic;
        C405DBGWBIAR05  : out    vl_logic;
        C405DBGWBIAR06  : out    vl_logic;
        C405DBGWBIAR07  : out    vl_logic;
        C405DBGWBIAR08  : out    vl_logic;
        C405DBGWBIAR09  : out    vl_logic;
        C405DBGWBIAR10  : out    vl_logic;
        C405DBGWBIAR11  : out    vl_logic;
        C405DBGWBIAR12  : out    vl_logic;
        C405DBGWBIAR13  : out    vl_logic;
        C405DBGWBIAR14  : out    vl_logic;
        C405DBGWBIAR15  : out    vl_logic;
        C405DBGWBIAR16  : out    vl_logic;
        C405DBGWBIAR17  : out    vl_logic;
        C405DBGWBIAR18  : out    vl_logic;
        C405DBGWBIAR19  : out    vl_logic;
        C405DBGWBIAR20  : out    vl_logic;
        C405DBGWBIAR21  : out    vl_logic;
        C405DBGWBIAR22  : out    vl_logic;
        C405DBGWBIAR23  : out    vl_logic;
        C405DBGWBIAR24  : out    vl_logic;
        C405DBGWBIAR25  : out    vl_logic;
        C405DBGWBIAR26  : out    vl_logic;
        C405DBGWBIAR27  : out    vl_logic;
        C405DBGWBIAR28  : out    vl_logic;
        C405DBGWBIAR29  : out    vl_logic;
        C405DCRABUS0    : out    vl_logic;
        C405DCRABUS1    : out    vl_logic;
        C405DCRABUS2    : out    vl_logic;
        C405DCRABUS3    : out    vl_logic;
        C405DCRABUS4    : out    vl_logic;
        C405DCRABUS5    : out    vl_logic;
        C405DCRABUS6    : out    vl_logic;
        C405DCRABUS7    : out    vl_logic;
        C405DCRABUS8    : out    vl_logic;
        C405DCRABUS9    : out    vl_logic;
        C405DCRDBUSOUT00: out    vl_logic;
        C405DCRDBUSOUT01: out    vl_logic;
        C405DCRDBUSOUT02: out    vl_logic;
        C405DCRDBUSOUT03: out    vl_logic;
        C405DCRDBUSOUT04: out    vl_logic;
        C405DCRDBUSOUT05: out    vl_logic;
        C405DCRDBUSOUT06: out    vl_logic;
        C405DCRDBUSOUT07: out    vl_logic;
        C405DCRDBUSOUT08: out    vl_logic;
        C405DCRDBUSOUT09: out    vl_logic;
        C405DCRDBUSOUT10: out    vl_logic;
        C405DCRDBUSOUT11: out    vl_logic;
        C405DCRDBUSOUT12: out    vl_logic;
        C405DCRDBUSOUT13: out    vl_logic;
        C405DCRDBUSOUT14: out    vl_logic;
        C405DCRDBUSOUT15: out    vl_logic;
        C405DCRDBUSOUT16: out    vl_logic;
        C405DCRDBUSOUT17: out    vl_logic;
        C405DCRDBUSOUT18: out    vl_logic;
        C405DCRDBUSOUT19: out    vl_logic;
        C405DCRDBUSOUT20: out    vl_logic;
        C405DCRDBUSOUT21: out    vl_logic;
        C405DCRDBUSOUT22: out    vl_logic;
        C405DCRDBUSOUT23: out    vl_logic;
        C405DCRDBUSOUT24: out    vl_logic;
        C405DCRDBUSOUT25: out    vl_logic;
        C405DCRDBUSOUT26: out    vl_logic;
        C405DCRDBUSOUT27: out    vl_logic;
        C405DCRDBUSOUT28: out    vl_logic;
        C405DCRDBUSOUT29: out    vl_logic;
        C405DCRDBUSOUT30: out    vl_logic;
        C405DCRDBUSOUT31: out    vl_logic;
        C405DCRREAD     : out    vl_logic;
        C405DCRWRITE    : out    vl_logic;
        C405DSOCMABORTOP: out    vl_logic;
        C405DSOCMABORTREQ: out    vl_logic;
        C405DSOCMABUS00 : out    vl_logic;
        C405DSOCMABUS01 : out    vl_logic;
        C405DSOCMABUS02 : out    vl_logic;
        C405DSOCMABUS03 : out    vl_logic;
        C405DSOCMABUS04 : out    vl_logic;
        C405DSOCMABUS05 : out    vl_logic;
        C405DSOCMABUS06 : out    vl_logic;
        C405DSOCMABUS07 : out    vl_logic;
        C405DSOCMABUS08 : out    vl_logic;
        C405DSOCMABUS09 : out    vl_logic;
        C405DSOCMABUS10 : out    vl_logic;
        C405DSOCMABUS11 : out    vl_logic;
        C405DSOCMABUS12 : out    vl_logic;
        C405DSOCMABUS13 : out    vl_logic;
        C405DSOCMABUS14 : out    vl_logic;
        C405DSOCMABUS15 : out    vl_logic;
        C405DSOCMABUS16 : out    vl_logic;
        C405DSOCMABUS17 : out    vl_logic;
        C405DSOCMABUS18 : out    vl_logic;
        C405DSOCMABUS19 : out    vl_logic;
        C405DSOCMABUS20 : out    vl_logic;
        C405DSOCMABUS21 : out    vl_logic;
        C405DSOCMABUS22 : out    vl_logic;
        C405DSOCMABUS23 : out    vl_logic;
        C405DSOCMABUS24 : out    vl_logic;
        C405DSOCMABUS25 : out    vl_logic;
        C405DSOCMABUS26 : out    vl_logic;
        C405DSOCMABUS27 : out    vl_logic;
        C405DSOCMABUS28 : out    vl_logic;
        C405DSOCMABUS29 : out    vl_logic;
        C405DSOCMBYTEEN0: out    vl_logic;
        C405DSOCMBYTEEN1: out    vl_logic;
        C405DSOCMBYTEEN2: out    vl_logic;
        C405DSOCMBYTEEN3: out    vl_logic;
        C405DSOCMCACHEABLE: out    vl_logic;
        C405DSOCMGUARDED: out    vl_logic;
        C405DSOCMLOADREQ: out    vl_logic;
        C405DSOCMSTOREREQ: out    vl_logic;
        C405DSOCMSTRINGMULTIPLE: out    vl_logic;
        C405DSOCMU0ATTR : out    vl_logic;
        C405DSOCMWAIT   : out    vl_logic;
        C405DSOCMWRDBUS00: out    vl_logic;
        C405DSOCMWRDBUS01: out    vl_logic;
        C405DSOCMWRDBUS02: out    vl_logic;
        C405DSOCMWRDBUS03: out    vl_logic;
        C405DSOCMWRDBUS04: out    vl_logic;
        C405DSOCMWRDBUS05: out    vl_logic;
        C405DSOCMWRDBUS06: out    vl_logic;
        C405DSOCMWRDBUS07: out    vl_logic;
        C405DSOCMWRDBUS08: out    vl_logic;
        C405DSOCMWRDBUS09: out    vl_logic;
        C405DSOCMWRDBUS10: out    vl_logic;
        C405DSOCMWRDBUS11: out    vl_logic;
        C405DSOCMWRDBUS12: out    vl_logic;
        C405DSOCMWRDBUS13: out    vl_logic;
        C405DSOCMWRDBUS14: out    vl_logic;
        C405DSOCMWRDBUS15: out    vl_logic;
        C405DSOCMWRDBUS16: out    vl_logic;
        C405DSOCMWRDBUS17: out    vl_logic;
        C405DSOCMWRDBUS18: out    vl_logic;
        C405DSOCMWRDBUS19: out    vl_logic;
        C405DSOCMWRDBUS20: out    vl_logic;
        C405DSOCMWRDBUS21: out    vl_logic;
        C405DSOCMWRDBUS22: out    vl_logic;
        C405DSOCMWRDBUS23: out    vl_logic;
        C405DSOCMWRDBUS24: out    vl_logic;
        C405DSOCMWRDBUS25: out    vl_logic;
        C405DSOCMWRDBUS26: out    vl_logic;
        C405DSOCMWRDBUS27: out    vl_logic;
        C405DSOCMWRDBUS28: out    vl_logic;
        C405DSOCMWRDBUS29: out    vl_logic;
        C405DSOCMWRDBUS30: out    vl_logic;
        C405DSOCMWRDBUS31: out    vl_logic;
        C405DSOCMXLATEVALID: out    vl_logic;
        C405ISOCMABORT  : out    vl_logic;
        C405ISOCMABUS00 : out    vl_logic;
        C405ISOCMABUS01 : out    vl_logic;
        C405ISOCMABUS02 : out    vl_logic;
        C405ISOCMABUS03 : out    vl_logic;
        C405ISOCMABUS04 : out    vl_logic;
        C405ISOCMABUS05 : out    vl_logic;
        C405ISOCMABUS06 : out    vl_logic;
        C405ISOCMABUS07 : out    vl_logic;
        C405ISOCMABUS08 : out    vl_logic;
        C405ISOCMABUS09 : out    vl_logic;
        C405ISOCMABUS10 : out    vl_logic;
        C405ISOCMABUS11 : out    vl_logic;
        C405ISOCMABUS12 : out    vl_logic;
        C405ISOCMABUS13 : out    vl_logic;
        C405ISOCMABUS14 : out    vl_logic;
        C405ISOCMABUS15 : out    vl_logic;
        C405ISOCMABUS16 : out    vl_logic;
        C405ISOCMABUS17 : out    vl_logic;
        C405ISOCMABUS18 : out    vl_logic;
        C405ISOCMABUS19 : out    vl_logic;
        C405ISOCMABUS20 : out    vl_logic;
        C405ISOCMABUS21 : out    vl_logic;
        C405ISOCMABUS22 : out    vl_logic;
        C405ISOCMABUS23 : out    vl_logic;
        C405ISOCMABUS24 : out    vl_logic;
        C405ISOCMABUS25 : out    vl_logic;
        C405ISOCMABUS26 : out    vl_logic;
        C405ISOCMABUS27 : out    vl_logic;
        C405ISOCMABUS28 : out    vl_logic;
        C405ISOCMABUS29 : out    vl_logic;
        C405ISOCMCACHEABLE: out    vl_logic;
        C405ISOCMCONTEXTSYNC: out    vl_logic;
        C405ISOCMICUREADY: out    vl_logic;
        C405ISOCMREQPENDING: out    vl_logic;
        C405ISOCMU0ATTR : out    vl_logic;
        C405ISOCMXLATEVALID: out    vl_logic;
        C405JTGCAPTUREDR: out    vl_logic;
        C405JTGEXTEST   : out    vl_logic;
        C405JTGPGMOUT   : out    vl_logic;
        C405JTGSHIFTDR  : out    vl_logic;
        C405JTGTDO      : out    vl_logic;
        C405JTGTDOEN    : out    vl_logic;
        C405JTGUPDATEDR : out    vl_logic;
        C405TESTDIAGABISTDONE: out    vl_logic;
        C405TESTSCANOUT0: out    vl_logic;
        C405TESTSCANOUT1: out    vl_logic;
        C405TESTSCANOUT2: out    vl_logic;
        C405TESTSCANOUT3: out    vl_logic;
        C405TESTSCANOUT4: out    vl_logic;
        C405TESTSCANOUT5: out    vl_logic;
        C405TESTSCANOUT6: out    vl_logic;
        C405TESTSCANOUT7: out    vl_logic;
        C405PLBDCUABORT : out    vl_logic;
        C405PLBDCUABUS00: out    vl_logic;
        C405PLBDCUABUS01: out    vl_logic;
        C405PLBDCUABUS02: out    vl_logic;
        C405PLBDCUABUS03: out    vl_logic;
        C405PLBDCUABUS04: out    vl_logic;
        C405PLBDCUABUS05: out    vl_logic;
        C405PLBDCUABUS06: out    vl_logic;
        C405PLBDCUABUS07: out    vl_logic;
        C405PLBDCUABUS08: out    vl_logic;
        C405PLBDCUABUS09: out    vl_logic;
        C405PLBDCUABUS10: out    vl_logic;
        C405PLBDCUABUS11: out    vl_logic;
        C405PLBDCUABUS12: out    vl_logic;
        C405PLBDCUABUS13: out    vl_logic;
        C405PLBDCUABUS14: out    vl_logic;
        C405PLBDCUABUS15: out    vl_logic;
        C405PLBDCUABUS16: out    vl_logic;
        C405PLBDCUABUS17: out    vl_logic;
        C405PLBDCUABUS18: out    vl_logic;
        C405PLBDCUABUS19: out    vl_logic;
        C405PLBDCUABUS20: out    vl_logic;
        C405PLBDCUABUS21: out    vl_logic;
        C405PLBDCUABUS22: out    vl_logic;
        C405PLBDCUABUS23: out    vl_logic;
        C405PLBDCUABUS24: out    vl_logic;
        C405PLBDCUABUS25: out    vl_logic;
        C405PLBDCUABUS26: out    vl_logic;
        C405PLBDCUABUS27: out    vl_logic;
        C405PLBDCUABUS28: out    vl_logic;
        C405PLBDCUABUS29: out    vl_logic;
        C405PLBDCUABUS30: out    vl_logic;
        C405PLBDCUABUS31: out    vl_logic;
        C405PLBDCUBE0   : out    vl_logic;
        C405PLBDCUBE1   : out    vl_logic;
        C405PLBDCUBE2   : out    vl_logic;
        C405PLBDCUBE3   : out    vl_logic;
        C405PLBDCUBE4   : out    vl_logic;
        C405PLBDCUBE5   : out    vl_logic;
        C405PLBDCUBE6   : out    vl_logic;
        C405PLBDCUBE7   : out    vl_logic;
        C405PLBDCUCACHEABLE: out    vl_logic;
        C405PLBDCUGUARDED: out    vl_logic;
        C405PLBDCUPRIORITY0: out    vl_logic;
        C405PLBDCUPRIORITY1: out    vl_logic;
        C405PLBDCUREQUEST: out    vl_logic;
        C405PLBDCURNW   : out    vl_logic;
        C405PLBDCUSIZE2 : out    vl_logic;
        C405PLBDCUU0ATTR: out    vl_logic;
        C405PLBDCUWRDBUS00: out    vl_logic;
        C405PLBDCUWRDBUS01: out    vl_logic;
        C405PLBDCUWRDBUS02: out    vl_logic;
        C405PLBDCUWRDBUS03: out    vl_logic;
        C405PLBDCUWRDBUS04: out    vl_logic;
        C405PLBDCUWRDBUS05: out    vl_logic;
        C405PLBDCUWRDBUS06: out    vl_logic;
        C405PLBDCUWRDBUS07: out    vl_logic;
        C405PLBDCUWRDBUS08: out    vl_logic;
        C405PLBDCUWRDBUS09: out    vl_logic;
        C405PLBDCUWRDBUS10: out    vl_logic;
        C405PLBDCUWRDBUS11: out    vl_logic;
        C405PLBDCUWRDBUS12: out    vl_logic;
        C405PLBDCUWRDBUS13: out    vl_logic;
        C405PLBDCUWRDBUS14: out    vl_logic;
        C405PLBDCUWRDBUS15: out    vl_logic;
        C405PLBDCUWRDBUS16: out    vl_logic;
        C405PLBDCUWRDBUS17: out    vl_logic;
        C405PLBDCUWRDBUS18: out    vl_logic;
        C405PLBDCUWRDBUS19: out    vl_logic;
        C405PLBDCUWRDBUS20: out    vl_logic;
        C405PLBDCUWRDBUS21: out    vl_logic;
        C405PLBDCUWRDBUS22: out    vl_logic;
        C405PLBDCUWRDBUS23: out    vl_logic;
        C405PLBDCUWRDBUS24: out    vl_logic;
        C405PLBDCUWRDBUS25: out    vl_logic;
        C405PLBDCUWRDBUS26: out    vl_logic;
        C405PLBDCUWRDBUS27: out    vl_logic;
        C405PLBDCUWRDBUS28: out    vl_logic;
        C405PLBDCUWRDBUS29: out    vl_logic;
        C405PLBDCUWRDBUS30: out    vl_logic;
        C405PLBDCUWRDBUS31: out    vl_logic;
        C405PLBDCUWRDBUS32: out    vl_logic;
        C405PLBDCUWRDBUS33: out    vl_logic;
        C405PLBDCUWRDBUS34: out    vl_logic;
        C405PLBDCUWRDBUS35: out    vl_logic;
        C405PLBDCUWRDBUS36: out    vl_logic;
        C405PLBDCUWRDBUS37: out    vl_logic;
        C405PLBDCUWRDBUS38: out    vl_logic;
        C405PLBDCUWRDBUS39: out    vl_logic;
        C405PLBDCUWRDBUS40: out    vl_logic;
        C405PLBDCUWRDBUS41: out    vl_logic;
        C405PLBDCUWRDBUS42: out    vl_logic;
        C405PLBDCUWRDBUS43: out    vl_logic;
        C405PLBDCUWRDBUS44: out    vl_logic;
        C405PLBDCUWRDBUS45: out    vl_logic;
        C405PLBDCUWRDBUS46: out    vl_logic;
        C405PLBDCUWRDBUS47: out    vl_logic;
        C405PLBDCUWRDBUS48: out    vl_logic;
        C405PLBDCUWRDBUS49: out    vl_logic;
        C405PLBDCUWRDBUS50: out    vl_logic;
        C405PLBDCUWRDBUS51: out    vl_logic;
        C405PLBDCUWRDBUS52: out    vl_logic;
        C405PLBDCUWRDBUS53: out    vl_logic;
        C405PLBDCUWRDBUS54: out    vl_logic;
        C405PLBDCUWRDBUS55: out    vl_logic;
        C405PLBDCUWRDBUS56: out    vl_logic;
        C405PLBDCUWRDBUS57: out    vl_logic;
        C405PLBDCUWRDBUS58: out    vl_logic;
        C405PLBDCUWRDBUS59: out    vl_logic;
        C405PLBDCUWRDBUS60: out    vl_logic;
        C405PLBDCUWRDBUS61: out    vl_logic;
        C405PLBDCUWRDBUS62: out    vl_logic;
        C405PLBDCUWRDBUS63: out    vl_logic;
        C405PLBDCUWRITETHRU: out    vl_logic;
        C405PLBICUABORT : out    vl_logic;
        C405PLBICUABUS00: out    vl_logic;
        C405PLBICUABUS01: out    vl_logic;
        C405PLBICUABUS02: out    vl_logic;
        C405PLBICUABUS03: out    vl_logic;
        C405PLBICUABUS04: out    vl_logic;
        C405PLBICUABUS05: out    vl_logic;
        C405PLBICUABUS06: out    vl_logic;
        C405PLBICUABUS07: out    vl_logic;
        C405PLBICUABUS08: out    vl_logic;
        C405PLBICUABUS09: out    vl_logic;
        C405PLBICUABUS10: out    vl_logic;
        C405PLBICUABUS11: out    vl_logic;
        C405PLBICUABUS12: out    vl_logic;
        C405PLBICUABUS13: out    vl_logic;
        C405PLBICUABUS14: out    vl_logic;
        C405PLBICUABUS15: out    vl_logic;
        C405PLBICUABUS16: out    vl_logic;
        C405PLBICUABUS17: out    vl_logic;
        C405PLBICUABUS18: out    vl_logic;
        C405PLBICUABUS19: out    vl_logic;
        C405PLBICUABUS20: out    vl_logic;
        C405PLBICUABUS21: out    vl_logic;
        C405PLBICUABUS22: out    vl_logic;
        C405PLBICUABUS23: out    vl_logic;
        C405PLBICUABUS24: out    vl_logic;
        C405PLBICUABUS25: out    vl_logic;
        C405PLBICUABUS26: out    vl_logic;
        C405PLBICUABUS27: out    vl_logic;
        C405PLBICUABUS28: out    vl_logic;
        C405PLBICUABUS29: out    vl_logic;
        C405PLBICUCACHEABLE: out    vl_logic;
        C405PLBICUPRIORITY0: out    vl_logic;
        C405PLBICUPRIORITY1: out    vl_logic;
        C405PLBICUREQUEST: out    vl_logic;
        C405PLBICUSIZE2 : out    vl_logic;
        C405PLBICUSIZE3 : out    vl_logic;
        C405PLBICUU0ATTR: out    vl_logic;
        C405RSTCHIPRESETREQ: out    vl_logic;
        C405RSTCORERESETREQ: out    vl_logic;
        C405RSTSYSTEMRESETREQ: out    vl_logic;
        C405TRCCYCLE    : out    vl_logic;
        C405TRCEVENEXECUTIONSTATUS0: out    vl_logic;
        C405TRCEVENEXECUTIONSTATUS1: out    vl_logic;
        C405TRCODDEXECUTIONSTATUS0: out    vl_logic;
        C405TRCODDEXECUTIONSTATUS1: out    vl_logic;
        C405TRCTRACESTATUS0: out    vl_logic;
        C405TRCTRACESTATUS1: out    vl_logic;
        C405TRCTRACESTATUS2: out    vl_logic;
        C405TRCTRACESTATUS3: out    vl_logic;
        C405TRCTRIGGEREVENTOUT: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE0: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE1: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE2: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE3: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE4: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE5: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE6: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE7: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE8: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE9: out    vl_logic;
        C405TRCTRIGGEREVENTTYPE10: out    vl_logic;
        C405XXXMACHINECHECK: out    vl_logic;
        APUC405DCDAPUOP : in     vl_logic;
        APUC405DCDCREN  : in     vl_logic;
        APUC405DCDFORCEALGN: in     vl_logic;
        APUC405DCDFORCEBESTEERING: in     vl_logic;
        APUC405DCDFPUOP : in     vl_logic;
        APUC405DCDGPRWRITE: in     vl_logic;
        APUC405DCDLDSTBYTE: in     vl_logic;
        APUC405DCDLDSTDW: in     vl_logic;
        APUC405DCDLDSTHW: in     vl_logic;
        APUC405DCDLDSTQW: in     vl_logic;
        APUC405DCDLDSTWD: in     vl_logic;
        APUC405DCDLOAD  : in     vl_logic;
        APUC405DCDPRIVOP: in     vl_logic;
        APUC405DCDRAEN  : in     vl_logic;
        APUC405DCDRBEN  : in     vl_logic;
        APUC405DCDSTORE : in     vl_logic;
        APUC405DCDTRAPBE: in     vl_logic;
        APUC405DCDTRAPLE: in     vl_logic;
        APUC405DCDUPDATE: in     vl_logic;
        APUC405DCDVALIDOP: in     vl_logic;
        APUC405DCDXERCAEN: in     vl_logic;
        APUC405DCDXEROVEN: in     vl_logic;
        APUC405EXCEPTION: in     vl_logic;
        APUC405EXEBLOCKINGMCO: in     vl_logic;
        APUC405EXEBUSY  : in     vl_logic;
        APUC405EXECR0   : in     vl_logic;
        APUC405EXECR1   : in     vl_logic;
        APUC405EXECR2   : in     vl_logic;
        APUC405EXECR3   : in     vl_logic;
        APUC405EXECRFIELD0: in     vl_logic;
        APUC405EXECRFIELD1: in     vl_logic;
        APUC405EXECRFIELD2: in     vl_logic;
        APUC405EXELDDEPEND: in     vl_logic;
        APUC405EXENONBLOCKINGMCO: in     vl_logic;
        APUC405EXERESULT00: in     vl_logic;
        APUC405EXERESULT01: in     vl_logic;
        APUC405EXERESULT02: in     vl_logic;
        APUC405EXERESULT03: in     vl_logic;
        APUC405EXERESULT04: in     vl_logic;
        APUC405EXERESULT05: in     vl_logic;
        APUC405EXERESULT06: in     vl_logic;
        APUC405EXERESULT07: in     vl_logic;
        APUC405EXERESULT08: in     vl_logic;
        APUC405EXERESULT09: in     vl_logic;
        APUC405EXERESULT10: in     vl_logic;
        APUC405EXERESULT11: in     vl_logic;
        APUC405EXERESULT12: in     vl_logic;
        APUC405EXERESULT13: in     vl_logic;
        APUC405EXERESULT14: in     vl_logic;
        APUC405EXERESULT15: in     vl_logic;
        APUC405EXERESULT16: in     vl_logic;
        APUC405EXERESULT17: in     vl_logic;
        APUC405EXERESULT18: in     vl_logic;
        APUC405EXERESULT19: in     vl_logic;
        APUC405EXERESULT20: in     vl_logic;
        APUC405EXERESULT21: in     vl_logic;
        APUC405EXERESULT22: in     vl_logic;
        APUC405EXERESULT23: in     vl_logic;
        APUC405EXERESULT24: in     vl_logic;
        APUC405EXERESULT25: in     vl_logic;
        APUC405EXERESULT26: in     vl_logic;
        APUC405EXERESULT27: in     vl_logic;
        APUC405EXERESULT28: in     vl_logic;
        APUC405EXERESULT29: in     vl_logic;
        APUC405EXERESULT30: in     vl_logic;
        APUC405EXERESULT31: in     vl_logic;
        APUC405EXEXERCA : in     vl_logic;
        APUC405EXEXEROV : in     vl_logic;
        APUC405FPUEXCEPTION: in     vl_logic;
        APUC405LWBLDDEPEND: in     vl_logic;
        APUC405SLEEPREQ : in     vl_logic;
        APUC405WBLDDEPEND: in     vl_logic;
        CPMC405CLOCK    : in     vl_logic;
        CPMC405CPUCLKENCCLK: in     vl_logic;
        CPMC405CORECLKINACTIVE: in     vl_logic;
        CPMC405JTAGCLKENCCLK: in     vl_logic;
        CPMC405PLBSAMPLECYCLE: in     vl_logic;
        CPMC405TIMERCLKENCCLK: in     vl_logic;
        CPMC405TIMERTICK: in     vl_logic;
        DBGC405DEBUGHALT: in     vl_logic;
        DBGC405EXTBUSHOLDACK: in     vl_logic;
        DBGC405UNCONDDEBUGEVENT: in     vl_logic;
        DCRC405ACK      : in     vl_logic;
        DCRC405DBUSIN00 : in     vl_logic;
        DCRC405DBUSIN01 : in     vl_logic;
        DCRC405DBUSIN02 : in     vl_logic;
        DCRC405DBUSIN03 : in     vl_logic;
        DCRC405DBUSIN04 : in     vl_logic;
        DCRC405DBUSIN05 : in     vl_logic;
        DCRC405DBUSIN06 : in     vl_logic;
        DCRC405DBUSIN07 : in     vl_logic;
        DCRC405DBUSIN08 : in     vl_logic;
        DCRC405DBUSIN09 : in     vl_logic;
        DCRC405DBUSIN10 : in     vl_logic;
        DCRC405DBUSIN11 : in     vl_logic;
        DCRC405DBUSIN12 : in     vl_logic;
        DCRC405DBUSIN13 : in     vl_logic;
        DCRC405DBUSIN14 : in     vl_logic;
        DCRC405DBUSIN15 : in     vl_logic;
        DCRC405DBUSIN16 : in     vl_logic;
        DCRC405DBUSIN17 : in     vl_logic;
        DCRC405DBUSIN18 : in     vl_logic;
        DCRC405DBUSIN19 : in     vl_logic;
        DCRC405DBUSIN20 : in     vl_logic;
        DCRC405DBUSIN21 : in     vl_logic;
        DCRC405DBUSIN22 : in     vl_logic;
        DCRC405DBUSIN23 : in     vl_logic;
        DCRC405DBUSIN24 : in     vl_logic;
        DCRC405DBUSIN25 : in     vl_logic;
        DCRC405DBUSIN26 : in     vl_logic;
        DCRC405DBUSIN27 : in     vl_logic;
        DCRC405DBUSIN28 : in     vl_logic;
        DCRC405DBUSIN29 : in     vl_logic;
        DCRC405DBUSIN30 : in     vl_logic;
        DCRC405DBUSIN31 : in     vl_logic;
        DSOCMC405COMPLETE: in     vl_logic;
        DSOCMC405DISOPERANDFWD: in     vl_logic;
        DSOCMC405HOLD   : in     vl_logic;
        DSOCMC405RDDBUS00: in     vl_logic;
        DSOCMC405RDDBUS01: in     vl_logic;
        DSOCMC405RDDBUS02: in     vl_logic;
        DSOCMC405RDDBUS03: in     vl_logic;
        DSOCMC405RDDBUS04: in     vl_logic;
        DSOCMC405RDDBUS05: in     vl_logic;
        DSOCMC405RDDBUS06: in     vl_logic;
        DSOCMC405RDDBUS07: in     vl_logic;
        DSOCMC405RDDBUS08: in     vl_logic;
        DSOCMC405RDDBUS09: in     vl_logic;
        DSOCMC405RDDBUS10: in     vl_logic;
        DSOCMC405RDDBUS11: in     vl_logic;
        DSOCMC405RDDBUS12: in     vl_logic;
        DSOCMC405RDDBUS13: in     vl_logic;
        DSOCMC405RDDBUS14: in     vl_logic;
        DSOCMC405RDDBUS15: in     vl_logic;
        DSOCMC405RDDBUS16: in     vl_logic;
        DSOCMC405RDDBUS17: in     vl_logic;
        DSOCMC405RDDBUS18: in     vl_logic;
        DSOCMC405RDDBUS19: in     vl_logic;
        DSOCMC405RDDBUS20: in     vl_logic;
        DSOCMC405RDDBUS21: in     vl_logic;
        DSOCMC405RDDBUS22: in     vl_logic;
        DSOCMC405RDDBUS23: in     vl_logic;
        DSOCMC405RDDBUS24: in     vl_logic;
        DSOCMC405RDDBUS25: in     vl_logic;
        DSOCMC405RDDBUS26: in     vl_logic;
        DSOCMC405RDDBUS27: in     vl_logic;
        DSOCMC405RDDBUS28: in     vl_logic;
        DSOCMC405RDDBUS29: in     vl_logic;
        DSOCMC405RDDBUS30: in     vl_logic;
        DSOCMC405RDDBUS31: in     vl_logic;
        EICC405CRITINPUTIRQ: in     vl_logic;
        EICC405EXTINPUTIRQ: in     vl_logic;
        ISOCMC405HOLD   : in     vl_logic;
        ISOCMC405RDDBUS00: in     vl_logic;
        ISOCMC405RDDBUS01: in     vl_logic;
        ISOCMC405RDDBUS02: in     vl_logic;
        ISOCMC405RDDBUS03: in     vl_logic;
        ISOCMC405RDDBUS04: in     vl_logic;
        ISOCMC405RDDBUS05: in     vl_logic;
        ISOCMC405RDDBUS06: in     vl_logic;
        ISOCMC405RDDBUS07: in     vl_logic;
        ISOCMC405RDDBUS08: in     vl_logic;
        ISOCMC405RDDBUS09: in     vl_logic;
        ISOCMC405RDDBUS10: in     vl_logic;
        ISOCMC405RDDBUS11: in     vl_logic;
        ISOCMC405RDDBUS12: in     vl_logic;
        ISOCMC405RDDBUS13: in     vl_logic;
        ISOCMC405RDDBUS14: in     vl_logic;
        ISOCMC405RDDBUS15: in     vl_logic;
        ISOCMC405RDDBUS16: in     vl_logic;
        ISOCMC405RDDBUS17: in     vl_logic;
        ISOCMC405RDDBUS18: in     vl_logic;
        ISOCMC405RDDBUS19: in     vl_logic;
        ISOCMC405RDDBUS20: in     vl_logic;
        ISOCMC405RDDBUS21: in     vl_logic;
        ISOCMC405RDDBUS22: in     vl_logic;
        ISOCMC405RDDBUS23: in     vl_logic;
        ISOCMC405RDDBUS24: in     vl_logic;
        ISOCMC405RDDBUS25: in     vl_logic;
        ISOCMC405RDDBUS26: in     vl_logic;
        ISOCMC405RDDBUS27: in     vl_logic;
        ISOCMC405RDDBUS28: in     vl_logic;
        ISOCMC405RDDBUS29: in     vl_logic;
        ISOCMC405RDDBUS30: in     vl_logic;
        ISOCMC405RDDBUS31: in     vl_logic;
        ISOCMC405RDDBUS32: in     vl_logic;
        ISOCMC405RDDBUS33: in     vl_logic;
        ISOCMC405RDDBUS34: in     vl_logic;
        ISOCMC405RDDBUS35: in     vl_logic;
        ISOCMC405RDDBUS36: in     vl_logic;
        ISOCMC405RDDBUS37: in     vl_logic;
        ISOCMC405RDDBUS38: in     vl_logic;
        ISOCMC405RDDBUS39: in     vl_logic;
        ISOCMC405RDDBUS40: in     vl_logic;
        ISOCMC405RDDBUS41: in     vl_logic;
        ISOCMC405RDDBUS42: in     vl_logic;
        ISOCMC405RDDBUS43: in     vl_logic;
        ISOCMC405RDDBUS44: in     vl_logic;
        ISOCMC405RDDBUS45: in     vl_logic;
        ISOCMC405RDDBUS46: in     vl_logic;
        ISOCMC405RDDBUS47: in     vl_logic;
        ISOCMC405RDDBUS48: in     vl_logic;
        ISOCMC405RDDBUS49: in     vl_logic;
        ISOCMC405RDDBUS50: in     vl_logic;
        ISOCMC405RDDBUS51: in     vl_logic;
        ISOCMC405RDDBUS52: in     vl_logic;
        ISOCMC405RDDBUS53: in     vl_logic;
        ISOCMC405RDDBUS54: in     vl_logic;
        ISOCMC405RDDBUS55: in     vl_logic;
        ISOCMC405RDDBUS56: in     vl_logic;
        ISOCMC405RDDBUS57: in     vl_logic;
        ISOCMC405RDDBUS58: in     vl_logic;
        ISOCMC405RDDBUS59: in     vl_logic;
        ISOCMC405RDDBUS60: in     vl_logic;
        ISOCMC405RDDBUS61: in     vl_logic;
        ISOCMC405RDDBUS62: in     vl_logic;
        ISOCMC405RDDBUS63: in     vl_logic;
        ISOCMC405RDDVALID0: in     vl_logic;
        ISOCMC405RDDVALID1: in     vl_logic;
        JTGC405BNDSCANTDO: in     vl_logic;
        JTGC405TCK      : in     vl_logic;
        JTGC405TDI      : in     vl_logic;
        JTGC405TMS      : in     vl_logic;
        JTGC405TRSTNEG  : in     vl_logic;
        TESTC405BISTCCLK: in     vl_logic;
        TESTC405SCANIN0 : in     vl_logic;
        TESTC405SCANIN1 : in     vl_logic;
        TESTC405SCANIN2 : in     vl_logic;
        TESTC405SCANIN3 : in     vl_logic;
        TESTC405SCANIN4 : in     vl_logic;
        TESTC405SCANIN5 : in     vl_logic;
        TESTC405SCANIN6 : in     vl_logic;
        TESTC405SCANIN7 : in     vl_logic;
        TESTC405SCANENABLE: in     vl_logic;
        TESTC405TESTMODE: in     vl_logic;
        TESTC405CNTLPOINT: in     vl_logic;
        TESTC405TESTM1  : in     vl_logic;
        TESTC405TESTM3  : in     vl_logic;
        PLBC405DCUADDRACK: in     vl_logic;
        PLBC405DCUBUSY  : in     vl_logic;
        PLBC405DCUERR   : in     vl_logic;
        PLBC405DCURDDACK: in     vl_logic;
        PLBC405DCURDDBUS00: in     vl_logic;
        PLBC405DCURDDBUS01: in     vl_logic;
        PLBC405DCURDDBUS02: in     vl_logic;
        PLBC405DCURDDBUS03: in     vl_logic;
        PLBC405DCURDDBUS04: in     vl_logic;
        PLBC405DCURDDBUS05: in     vl_logic;
        PLBC405DCURDDBUS06: in     vl_logic;
        PLBC405DCURDDBUS07: in     vl_logic;
        PLBC405DCURDDBUS08: in     vl_logic;
        PLBC405DCURDDBUS09: in     vl_logic;
        PLBC405DCURDDBUS10: in     vl_logic;
        PLBC405DCURDDBUS11: in     vl_logic;
        PLBC405DCURDDBUS12: in     vl_logic;
        PLBC405DCURDDBUS13: in     vl_logic;
        PLBC405DCURDDBUS14: in     vl_logic;
        PLBC405DCURDDBUS15: in     vl_logic;
        PLBC405DCURDDBUS16: in     vl_logic;
        PLBC405DCURDDBUS17: in     vl_logic;
        PLBC405DCURDDBUS18: in     vl_logic;
        PLBC405DCURDDBUS19: in     vl_logic;
        PLBC405DCURDDBUS20: in     vl_logic;
        PLBC405DCURDDBUS21: in     vl_logic;
        PLBC405DCURDDBUS22: in     vl_logic;
        PLBC405DCURDDBUS23: in     vl_logic;
        PLBC405DCURDDBUS24: in     vl_logic;
        PLBC405DCURDDBUS25: in     vl_logic;
        PLBC405DCURDDBUS26: in     vl_logic;
        PLBC405DCURDDBUS27: in     vl_logic;
        PLBC405DCURDDBUS28: in     vl_logic;
        PLBC405DCURDDBUS29: in     vl_logic;
        PLBC405DCURDDBUS30: in     vl_logic;
        PLBC405DCURDDBUS31: in     vl_logic;
        PLBC405DCURDDBUS32: in     vl_logic;
        PLBC405DCURDDBUS33: in     vl_logic;
        PLBC405DCURDDBUS34: in     vl_logic;
        PLBC405DCURDDBUS35: in     vl_logic;
        PLBC405DCURDDBUS36: in     vl_logic;
        PLBC405DCURDDBUS37: in     vl_logic;
        PLBC405DCURDDBUS38: in     vl_logic;
        PLBC405DCURDDBUS39: in     vl_logic;
        PLBC405DCURDDBUS40: in     vl_logic;
        PLBC405DCURDDBUS41: in     vl_logic;
        PLBC405DCURDDBUS42: in     vl_logic;
        PLBC405DCURDDBUS43: in     vl_logic;
        PLBC405DCURDDBUS44: in     vl_logic;
        PLBC405DCURDDBUS45: in     vl_logic;
        PLBC405DCURDDBUS46: in     vl_logic;
        PLBC405DCURDDBUS47: in     vl_logic;
        PLBC405DCURDDBUS48: in     vl_logic;
        PLBC405DCURDDBUS49: in     vl_logic;
        PLBC405DCURDDBUS50: in     vl_logic;
        PLBC405DCURDDBUS51: in     vl_logic;
        PLBC405DCURDDBUS52: in     vl_logic;
        PLBC405DCURDDBUS53: in     vl_logic;
        PLBC405DCURDDBUS54: in     vl_logic;
        PLBC405DCURDDBUS55: in     vl_logic;
        PLBC405DCURDDBUS56: in     vl_logic;
        PLBC405DCURDDBUS57: in     vl_logic;
        PLBC405DCURDDBUS58: in     vl_logic;
        PLBC405DCURDDBUS59: in     vl_logic;
        PLBC405DCURDDBUS60: in     vl_logic;
        PLBC405DCURDDBUS61: in     vl_logic;
        PLBC405DCURDDBUS62: in     vl_logic;
        PLBC405DCURDDBUS63: in     vl_logic;
        PLBC405DCURDWDADDR1: in     vl_logic;
        PLBC405DCURDWDADDR2: in     vl_logic;
        PLBC405DCURDWDADDR3: in     vl_logic;
        PLBC405DCUSSIZE1: in     vl_logic;
        PLBC405DCUWRDACK: in     vl_logic;
        PLBC405ICUADDRACK: in     vl_logic;
        PLBC405ICUBUSY  : in     vl_logic;
        PLBC405ICUERR   : in     vl_logic;
        PLBC405ICURDDACK: in     vl_logic;
        PLBC405ICURDDBUS00: in     vl_logic;
        PLBC405ICURDDBUS01: in     vl_logic;
        PLBC405ICURDDBUS02: in     vl_logic;
        PLBC405ICURDDBUS03: in     vl_logic;
        PLBC405ICURDDBUS04: in     vl_logic;
        PLBC405ICURDDBUS05: in     vl_logic;
        PLBC405ICURDDBUS06: in     vl_logic;
        PLBC405ICURDDBUS07: in     vl_logic;
        PLBC405ICURDDBUS08: in     vl_logic;
        PLBC405ICURDDBUS09: in     vl_logic;
        PLBC405ICURDDBUS10: in     vl_logic;
        PLBC405ICURDDBUS11: in     vl_logic;
        PLBC405ICURDDBUS12: in     vl_logic;
        PLBC405ICURDDBUS13: in     vl_logic;
        PLBC405ICURDDBUS14: in     vl_logic;
        PLBC405ICURDDBUS15: in     vl_logic;
        PLBC405ICURDDBUS16: in     vl_logic;
        PLBC405ICURDDBUS17: in     vl_logic;
        PLBC405ICURDDBUS18: in     vl_logic;
        PLBC405ICURDDBUS19: in     vl_logic;
        PLBC405ICURDDBUS20: in     vl_logic;
        PLBC405ICURDDBUS21: in     vl_logic;
        PLBC405ICURDDBUS22: in     vl_logic;
        PLBC405ICURDDBUS23: in     vl_logic;
        PLBC405ICURDDBUS24: in     vl_logic;
        PLBC405ICURDDBUS25: in     vl_logic;
        PLBC405ICURDDBUS26: in     vl_logic;
        PLBC405ICURDDBUS27: in     vl_logic;
        PLBC405ICURDDBUS28: in     vl_logic;
        PLBC405ICURDDBUS29: in     vl_logic;
        PLBC405ICURDDBUS30: in     vl_logic;
        PLBC405ICURDDBUS31: in     vl_logic;
        PLBC405ICURDDBUS32: in     vl_logic;
        PLBC405ICURDDBUS33: in     vl_logic;
        PLBC405ICURDDBUS34: in     vl_logic;
        PLBC405ICURDDBUS35: in     vl_logic;
        PLBC405ICURDDBUS36: in     vl_logic;
        PLBC405ICURDDBUS37: in     vl_logic;
        PLBC405ICURDDBUS38: in     vl_logic;
        PLBC405ICURDDBUS39: in     vl_logic;
        PLBC405ICURDDBUS40: in     vl_logic;
        PLBC405ICURDDBUS41: in     vl_logic;
        PLBC405ICURDDBUS42: in     vl_logic;
        PLBC405ICURDDBUS43: in     vl_logic;
        PLBC405ICURDDBUS44: in     vl_logic;
        PLBC405ICURDDBUS45: in     vl_logic;
        PLBC405ICURDDBUS46: in     vl_logic;
        PLBC405ICURDDBUS47: in     vl_logic;
        PLBC405ICURDDBUS48: in     vl_logic;
        PLBC405ICURDDBUS49: in     vl_logic;
        PLBC405ICURDDBUS50: in     vl_logic;
        PLBC405ICURDDBUS51: in     vl_logic;
        PLBC405ICURDDBUS52: in     vl_logic;
        PLBC405ICURDDBUS53: in     vl_logic;
        PLBC405ICURDDBUS54: in     vl_logic;
        PLBC405ICURDDBUS55: in     vl_logic;
        PLBC405ICURDDBUS56: in     vl_logic;
        PLBC405ICURDDBUS57: in     vl_logic;
        PLBC405ICURDDBUS58: in     vl_logic;
        PLBC405ICURDDBUS59: in     vl_logic;
        PLBC405ICURDDBUS60: in     vl_logic;
        PLBC405ICURDDBUS61: in     vl_logic;
        PLBC405ICURDDBUS62: in     vl_logic;
        PLBC405ICURDDBUS63: in     vl_logic;
        PLBC405ICURDWDADDR1: in     vl_logic;
        PLBC405ICURDWDADDR2: in     vl_logic;
        PLBC405ICURDWDADDR3: in     vl_logic;
        PLBC405ICUSSIZE1: in     vl_logic;
        RSTC405RESETCHIP: in     vl_logic;
        RSTC405RESETCORE: in     vl_logic;
        RSTC405RESETSYSTEM: in     vl_logic;
        TIEC405APUDIVEN : in     vl_logic;
        TIEC405APUPRESENT: in     vl_logic;
        TIEC405DETERMINISTICMULT: in     vl_logic;
        TIEC405DISOPERANDFWD: in     vl_logic;
        TIEC405MMUEN    : in     vl_logic;
        TIEC405PVR00    : in     vl_logic;
        TIEC405PVR01    : in     vl_logic;
        TIEC405PVR02    : in     vl_logic;
        TIEC405PVR03    : in     vl_logic;
        TIEC405PVR04    : in     vl_logic;
        TIEC405PVR05    : in     vl_logic;
        TIEC405PVR06    : in     vl_logic;
        TIEC405PVR07    : in     vl_logic;
        TIEC405PVR08    : in     vl_logic;
        TIEC405PVR09    : in     vl_logic;
        TIEC405PVR10    : in     vl_logic;
        TIEC405PVR11    : in     vl_logic;
        TIEC405PVR12    : in     vl_logic;
        TIEC405PVR13    : in     vl_logic;
        TIEC405PVR14    : in     vl_logic;
        TIEC405PVR15    : in     vl_logic;
        TIEC405PVR16    : in     vl_logic;
        TIEC405PVR17    : in     vl_logic;
        TIEC405PVR18    : in     vl_logic;
        TIEC405PVR19    : in     vl_logic;
        TIEC405PVR20    : in     vl_logic;
        TIEC405PVR21    : in     vl_logic;
        TIEC405PVR22    : in     vl_logic;
        TIEC405PVR23    : in     vl_logic;
        TIEC405PVR24    : in     vl_logic;
        TIEC405PVR25    : in     vl_logic;
        TIEC405PVR26    : in     vl_logic;
        TIEC405PVR27    : in     vl_logic;
        TIEC405PVR28    : in     vl_logic;
        TIEC405PVR29    : in     vl_logic;
        TIEC405PVR30    : in     vl_logic;
        TIEC405PVR31    : in     vl_logic;
        TRCC405TRACEDISABLE: in     vl_logic;
        TRCC405TRIGGEREVENTIN: in     vl_logic;
        C405BISTPEPSPF00: out    vl_logic;
        C405BISTPEPSPF01: out    vl_logic;
        C405BISTPEPSPF02: out    vl_logic;
        TESTC405CE0EVS  : in     vl_logic;
        TESTC405BISTCE0STCLK: in     vl_logic;
        TESTC405BISTCE1ENABLE: in     vl_logic;
        TESTC405BISTCE1MODE: in     vl_logic;
        CPMC405PLBSYNCCLOCK: in     vl_logic;
        CPMC405SYNCBYPASS: in     vl_logic;
        TIEC405CLOCKENABLE: in     vl_logic;
        TIEC405DUTYENABLE: in     vl_logic;
        CPMC405PLBSAMPLECYCLEALT: in     vl_logic;
        BISTC405DCUBISTDEBUGSI00: in     vl_logic;
        BISTC405DCUBISTDEBUGSI01: in     vl_logic;
        BISTC405DCUBISTDEBUGSI02: in     vl_logic;
        BISTC405DCUBISTDEBUGSI03: in     vl_logic;
        C405BISTDCUBISTDEBUGSO00: out    vl_logic;
        C405BISTDCUBISTDEBUGSO01: out    vl_logic;
        C405BISTDCUBISTDEBUGSO02: out    vl_logic;
        C405BISTDCUBISTDEBUGSO03: out    vl_logic;
        BISTC405DCUBISTDEBUGEN00: in     vl_logic;
        BISTC405DCUBISTDEBUGEN01: in     vl_logic;
        BISTC405DCUBISTDEBUGEN02: in     vl_logic;
        BISTC405DCUBISTDEBUGEN03: in     vl_logic;
        BISTC405DCUBISTMODEREGIN00: in     vl_logic;
        BISTC405DCUBISTMODEREGIN01: in     vl_logic;
        BISTC405DCUBISTMODEREGIN02: in     vl_logic;
        BISTC405DCUBISTMODEREGIN03: in     vl_logic;
        BISTC405DCUBISTMODEREGIN04: in     vl_logic;
        BISTC405DCUBISTMODEREGIN05: in     vl_logic;
        BISTC405DCUBISTMODEREGIN06: in     vl_logic;
        BISTC405DCUBISTMODEREGIN07: in     vl_logic;
        BISTC405DCUBISTMODEREGIN08: in     vl_logic;
        BISTC405DCUBISTMODEREGIN09: in     vl_logic;
        BISTC405DCUBISTMODEREGIN10: in     vl_logic;
        BISTC405DCUBISTMODEREGIN11: in     vl_logic;
        BISTC405DCUBISTMODEREGIN12: in     vl_logic;
        BISTC405DCUBISTMODEREGIN13: in     vl_logic;
        BISTC405DCUBISTMODEREGIN14: in     vl_logic;
        BISTC405DCUBISTMODEREGIN15: in     vl_logic;
        BISTC405DCUBISTMODEREGIN16: in     vl_logic;
        BISTC405DCUBISTMODEREGIN17: in     vl_logic;
        BISTC405DCUBISTMODEREGIN18: in     vl_logic;
        C405BISTDCUBISTMODEREGOUT00: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT01: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT02: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT03: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT04: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT05: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT06: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT07: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT08: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT09: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT10: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT11: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT12: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT13: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT14: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT15: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT16: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT17: out    vl_logic;
        C405BISTDCUBISTMODEREGOUT18: out    vl_logic;
        BISTC405DCUBISTMODEREGSI: in     vl_logic;
        C405BISTDCUBISTMODEREGSO: out    vl_logic;
        BISTC405DCUBISTSHIFTDR: in     vl_logic;
        BISTC405DCUBISTMBRUN: in     vl_logic;
        BISTC405DCUBISTPARALLELDR: in     vl_logic;
        BISTC405ICUBISTDEBUGSI00: in     vl_logic;
        BISTC405ICUBISTDEBUGSI01: in     vl_logic;
        BISTC405ICUBISTDEBUGSI02: in     vl_logic;
        BISTC405ICUBISTDEBUGSI03: in     vl_logic;
        C405BISTICUBISTDEBUGSO00: out    vl_logic;
        C405BISTICUBISTDEBUGSO01: out    vl_logic;
        C405BISTICUBISTDEBUGSO02: out    vl_logic;
        C405BISTICUBISTDEBUGSO03: out    vl_logic;
        BISTC405ICUBISTDEBUGEN00: in     vl_logic;
        BISTC405ICUBISTDEBUGEN01: in     vl_logic;
        BISTC405ICUBISTDEBUGEN02: in     vl_logic;
        BISTC405ICUBISTDEBUGEN03: in     vl_logic;
        BISTC405ICUBISTMODEREGIN00: in     vl_logic;
        BISTC405ICUBISTMODEREGIN01: in     vl_logic;
        BISTC405ICUBISTMODEREGIN02: in     vl_logic;
        BISTC405ICUBISTMODEREGIN03: in     vl_logic;
        BISTC405ICUBISTMODEREGIN04: in     vl_logic;
        BISTC405ICUBISTMODEREGIN05: in     vl_logic;
        BISTC405ICUBISTMODEREGIN06: in     vl_logic;
        BISTC405ICUBISTMODEREGIN07: in     vl_logic;
        BISTC405ICUBISTMODEREGIN08: in     vl_logic;
        BISTC405ICUBISTMODEREGIN09: in     vl_logic;
        BISTC405ICUBISTMODEREGIN10: in     vl_logic;
        BISTC405ICUBISTMODEREGIN11: in     vl_logic;
        BISTC405ICUBISTMODEREGIN12: in     vl_logic;
        BISTC405ICUBISTMODEREGIN13: in     vl_logic;
        BISTC405ICUBISTMODEREGIN14: in     vl_logic;
        BISTC405ICUBISTMODEREGIN15: in     vl_logic;
        BISTC405ICUBISTMODEREGIN16: in     vl_logic;
        BISTC405ICUBISTMODEREGIN17: in     vl_logic;
        BISTC405ICUBISTMODEREGIN18: in     vl_logic;
        C405BISTICUBISTMODEREGOUT00: out    vl_logic;
        C405BISTICUBISTMODEREGOUT01: out    vl_logic;
        C405BISTICUBISTMODEREGOUT02: out    vl_logic;
        C405BISTICUBISTMODEREGOUT03: out    vl_logic;
        C405BISTICUBISTMODEREGOUT04: out    vl_logic;
        C405BISTICUBISTMODEREGOUT05: out    vl_logic;
        C405BISTICUBISTMODEREGOUT06: out    vl_logic;
        C405BISTICUBISTMODEREGOUT07: out    vl_logic;
        C405BISTICUBISTMODEREGOUT08: out    vl_logic;
        C405BISTICUBISTMODEREGOUT09: out    vl_logic;
        C405BISTICUBISTMODEREGOUT10: out    vl_logic;
        C405BISTICUBISTMODEREGOUT11: out    vl_logic;
        C405BISTICUBISTMODEREGOUT12: out    vl_logic;
        C405BISTICUBISTMODEREGOUT13: out    vl_logic;
        C405BISTICUBISTMODEREGOUT14: out    vl_logic;
        C405BISTICUBISTMODEREGOUT15: out    vl_logic;
        C405BISTICUBISTMODEREGOUT16: out    vl_logic;
        C405BISTICUBISTMODEREGOUT17: out    vl_logic;
        C405BISTICUBISTMODEREGOUT18: out    vl_logic;
        BISTC405ICUBISTMODEREGSI: in     vl_logic;
        C405BISTICUBISTMODEREGSO: out    vl_logic;
        BISTC405ICUBISTSHIFTDR: in     vl_logic;
        BISTC405ICUBISTMBRUN: in     vl_logic;
        BISTC405ICUBISTPARALLELDR: in     vl_logic
    );
end PPC405F5V1;
