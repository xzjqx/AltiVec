library verilog;
use verilog.vl_types.all;
entity p405s_DTLB is
    port(
        CAR_Endian      : out    vl_logic;
        CAR_U0Attr      : out    vl_logic;
        CAR_XltValid    : out    vl_logic;
        CAR_cacheable   : out    vl_logic;
        CAR_guarded     : out    vl_logic;
        CAR_writethru   : out    vl_logic;
        DTLB_I          : out    vl_logic;
        DTLB_U0         : out    vl_logic;
        DTLB_W          : out    vl_logic;
        DTLB_WR         : out    vl_logic;
        DTLB_zonePR     : out    vl_logic_vector(0 to 1);
        MMU_apuWbEndian : out    vl_logic;
        MMU_rdarDsRAL2  : out    vl_logic_vector(0 to 29);
        dsRA            : out    vl_logic_vector(0 to 21);
        dtlbMiss        : out    vl_logic;
        isDsCacheableL2 : out    vl_logic;
        isDsEndianL2    : out    vl_logic;
        isDsU0AttrL2    : out    vl_logic;
        isDsXltValidL2  : out    vl_logic;
        CAR_mmuAttr_E1  : in     vl_logic;
        CAR_mmuAttr_E2  : in     vl_logic;
        CB              : in     vl_logic;
        DSize           : in     vl_logic_vector(0 to 6);
        E               : in     vl_logic;
        EXE_dsEaCP_NEG  : in     vl_logic_vector(0 to 7);
        EXE_eaARegBuf   : in     vl_logic_vector(0 to 21);
        EXE_eaBRegBuf   : in     vl_logic_vector(0 to 21);
        G               : in     vl_logic;
        I               : in     vl_logic;
        ICU_mmuRdarE2   : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        MMU_dsRA        : in     vl_logic_vector(22 to 29);
        RPN             : in     vl_logic_vector(0 to 21);
        U0              : in     vl_logic;
        W               : in     vl_logic;
        WR              : in     vl_logic;
        bypassRPN       : in     vl_logic_vector(0 to 21);
        dsAddr          : in     vl_logic_vector(0 to 2);
        dsEA_NEG        : in     vl_logic_vector(0 to 21);
        dsEPN           : in     vl_logic_vector(0 to 21);
        dsEReal_N       : in     vl_logic;
        dsGReal_N       : in     vl_logic;
        dsIReal_N       : in     vl_logic;
        dsInvalidate    : in     vl_logic;
        dsStateA        : in     vl_logic;
        dsStateD        : in     vl_logic;
        dsU0Real_N      : in     vl_logic;
        dsXltValid      : in     vl_logic;
        dsrdNotWrt      : in     vl_logic;
        isDsIReal_N     : in     vl_logic;
        msrDR           : in     vl_logic;
        wtReqReal_N     : in     vl_logic;
        zonePR          : in     vl_logic_vector(0 to 1)
    );
end p405s_DTLB;
