library verilog;
use verilog.vl_types.all;
entity p405s_pcl_top is
    port(
        PCL_LpEqSp      : out    vl_logic;
        PCL_Rbit        : out    vl_logic;
        PCL_aPortRregBypass: out    vl_logic;
        PCL_aRegE2      : out    vl_logic;
        PCL_aRegForEaE2 : out    vl_logic;
        PCL_abRegE1     : out    vl_logic;
        PCL_addFour     : out    vl_logic;
        PCL_apuDcdHold  : out    vl_logic;
        PCL_apuExeFlush : out    vl_logic;
        PCL_apuExeHold  : out    vl_logic;
        PCL_apuExeWdCnt : out    vl_logic_vector(0 to 1);
        PCL_apuLwbLoadDV: out    vl_logic;
        PCL_apuTrcLoadEn: out    vl_logic;
        PCL_apuWbHold   : out    vl_logic;
        PCL_bPortLitGenSel: out    vl_logic;
        PCL_bPortRregBypass: out    vl_logic;
        PCL_bRegE2      : out    vl_logic;
        PCL_bRegForEaE2 : out    vl_logic;
        PCL_blkFlush    : out    vl_logic;
        PCL_blkFlushForVct: out    vl_logic_vector(0 to 2);
        PCL_dIcmpForStep: out    vl_logic;
        PCL_dIcmpForStuff: out    vl_logic;
        PCL_dIcmpForWbFlushQDlydL2: out    vl_logic;
        PCL_dRegBypassMuxSel: out    vl_logic;
        PCL_dRegE1      : out    vl_logic;
        PCL_dbgSprDcds  : out    vl_logic_vector(0 to 3);
        PCL_dcdApAddr   : out    vl_logic_vector(0 to 9);
        PCL_dcdAregLoadUse: out    vl_logic;
        PCL_dcdBpAddr   : out    vl_logic_vector(0 to 9);
        PCL_dcdBregLoadUse: out    vl_logic;
        PCL_dcdHoldForIfb: out    vl_logic_vector(0 to 2);
        PCL_dcdHotCIn   : out    vl_logic;
        PCL_dcdImmd     : out    vl_logic_vector(11 to 31);
        PCL_dcdLitCntl  : out    vl_logic_vector(0 to 4);
        PCL_dcdMdSelQ   : out    vl_logic;
        PCL_dcdMrSelQ   : out    vl_logic;
        PCL_dcdSpAddr   : out    vl_logic_vector(0 to 9);
        PCL_dcdSregLoadUse: out    vl_logic;
        PCL_dcdSrmBpSel : out    vl_logic_vector(0 to 2);
        PCL_dcdXerCa    : out    vl_logic;
        PCL_dcuByteEn   : out    vl_logic_vector(0 to 3);
        PCL_dcuOp       : out    vl_logic_vector(0 to 11);
        PCL_dcuOp_early : out    vl_logic_vector(0 to 2);
        PCL_diagBus     : out    vl_logic_vector(0 to 9);
        PCL_dofDRegE1   : out    vl_logic;
        PCL_dofDRegMuxSel: out    vl_logic_vector(0 to 1);
        PCL_dsMmuOp     : out    vl_logic_vector(0 to 3);
        PCL_dsOcmByteEn : out    vl_logic_vector(0 to 3);
        PCL_dvcByteEnL2 : out    vl_logic_vector(0 to 3);
        PCL_dvcCmpEn    : out    vl_logic;
        PCL_exe2AccRegMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exe2ClearOrFlush: out    vl_logic;
        PCL_exe2DataE1  : out    vl_logic;
        PCL_exe2DataE2  : out    vl_logic;
        PCL_exe2Full    : out    vl_logic;
        PCL_exe2Hold    : out    vl_logic;
        PCL_exe2IarE1   : out    vl_logic;
        PCL_exe2IarE2   : out    vl_logic;
        PCL_exe2MacEn   : out    vl_logic;
        PCL_exe2MacOrMultEnForMS: out    vl_logic_vector(0 to 1);
        PCL_exe2MacOrMultEn_NEG: out    vl_logic_vector(0 to 1);
        PCL_exe2MacSat  : out    vl_logic;
        PCL_exe2MultEn  : out    vl_logic;
        PCL_exe2MultHiWd: out    vl_logic;
        PCL_exe2NegMac  : out    vl_logic;
        PCL_exe2SignedOp: out    vl_logic;
        PCL_exe2XerOvEn : out    vl_logic;
        PCL_exeAbort    : out    vl_logic;
        PCL_exeAddEn    : out    vl_logic;
        PCL_exeAddSgndOp_NEG: out    vl_logic_vector(0 to 1);
        PCL_exeAdmCntl  : out    vl_logic_vector(0 to 3);
        PCL_exeApuOp    : out    vl_logic;
        PCL_exeApuValidOp: out    vl_logic;
        PCL_exeAregLoadUse: out    vl_logic;
        PCL_exeBregLoadUse: out    vl_logic;
        PCL_exeCmplmntA : out    vl_logic;
        PCL_exeCmplmntA_NEG: out    vl_logic;
        PCL_exeCpuOp    : out    vl_logic;
        PCL_exeDbgLdOp  : out    vl_logic;
        PCL_exeDbgRdOp  : out    vl_logic;
        PCL_exeDbgStOp  : out    vl_logic;
        PCL_exeDbgWrOp  : out    vl_logic;
        PCL_exeDivEn    : out    vl_logic;
        PCL_exeDivEnForLSSD: out    vl_logic;
        PCL_exeDivEnForMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exeDivEn_NEG: out    vl_logic;
        PCL_exeDivSgndOp: out    vl_logic;
        PCL_exeDvcHold  : out    vl_logic;
        PCL_exeEaCalc   : out    vl_logic;
        PCL_exeEaQwEn   : out    vl_logic_vector(0 to 3);
        PCL_exeFpuOp    : out    vl_logic;
        PCL_exeFull     : out    vl_logic;
        PCL_exeHoldForCr: out    vl_logic;
        PCL_exeIarHold  : out    vl_logic;
        PCL_exeLdNotSt  : out    vl_logic;
        PCL_exeLoadUseHold: out    vl_logic;
        PCL_exeLogicalCntl: out    vl_logic_vector(0 to 7);
        PCL_exeLogicalUnitEnForLSSD: out    vl_logic;
        PCL_exeLogicalUnitEn_NEG: out    vl_logic;
        PCL_exeMacEn    : out    vl_logic;
        PCL_exeMacOrMultEn_NEG: out    vl_logic;
        PCL_exeMultEn   : out    vl_logic;
        PCL_exeMultEnForMuxSel: out    vl_logic_vector(0 to 1);
        PCL_exeMultEn_NEG: out    vl_logic_vector(0 to 1);
        PCL_exeNegMac   : out    vl_logic;
        PCL_exePrivOp   : out    vl_logic;
        PCL_exeRaEn     : out    vl_logic_vector(0 to 3);
        PCL_exeRbEn     : out    vl_logic_vector(0 to 3);
        PCL_exeSprDataEn_NEG: out    vl_logic;
        PCL_exeSprDcds  : out    vl_logic_vector(0 to 4);
        PCL_exeSprUnitEn_NEG: out    vl_logic;
        PCL_exeSregLoadUse: out    vl_logic;
        PCL_exeSrmBpSel : out    vl_logic_vector(0 to 2);
        PCL_exeSrmCntl  : out    vl_logic_vector(0 to 3);
        PCL_exeSrmUnitEnForLSSD: out    vl_logic;
        PCL_exeSrmUnitEn_NEG: out    vl_logic;
        PCL_exeStorageOp: out    vl_logic;
        PCL_exeStringMultiple: out    vl_logic;
        PCL_exeTlbOp    : out    vl_logic;
        PCL_exeTrap     : out    vl_logic;
        PCL_exeTrapCond : out    vl_logic_vector(0 to 4);
        PCL_exeWrExtEn  : out    vl_logic;
        PCL_exeWrtee    : out    vl_logic;
        PCL_exeXerCaEn  : out    vl_logic;
        PCL_exeXerOvEn  : out    vl_logic;
        PCL_gateZeroToAreg: out    vl_logic;
        PCL_gateZeroToSreg: out    vl_logic;
        PCL_holdCIn     : out    vl_logic;
        PCL_holdMdMr    : out    vl_logic;
        PCL_icuOp       : out    vl_logic_vector(0 to 3);
        PCL_icuSprDcds  : out    vl_logic_vector(0 to 2);
        PCL_ifbSprHold  : out    vl_logic;
        PCL_jtgSprDcd   : out    vl_logic;
        PCL_ldAdjE1     : out    vl_logic;
        PCL_ldAdjE2     : out    vl_logic_vector(1 to 3);
        PCL_ldAdjMuxSel : out    vl_logic_vector(0 to 1);
        PCL_ldFillBypassMuxSel: out    vl_logic_vector(0 to 5);
        PCL_ldMuxSel    : out    vl_logic_vector(0 to 7);
        PCL_ldSteerMuxSel: out    vl_logic_vector(0 to 7);
        PCL_lwbLpAddr   : out    vl_logic_vector(0 to 4);
        PCL_lwbLpEqdcdApAddr: out    vl_logic;
        PCL_lwbLpEqdcdBpAddr: out    vl_logic;
        PCL_lwbLpWrEn   : out    vl_logic;
        PCL_mfDCR       : out    vl_logic;
        PCL_mfDCRL2     : out    vl_logic;
        PCL_mfSPR       : out    vl_logic;
        PCL_mmuExeAbort : out    vl_logic;
        PCL_mmuIcuSprHold: out    vl_logic;
        PCL_mmuSprDcd   : out    vl_logic_vector(0 to 8);
        PCL_mtDCR       : out    vl_logic;
        PCL_mtSPR       : out    vl_logic;
        PCL_ocmAbortReq : out    vl_logic;
        PCL_resultMuxSel: out    vl_logic;
        PCL_resultRegE1 : out    vl_logic;
        PCL_resultRegE2 : out    vl_logic;
        PCL_sPortRregBypass: out    vl_logic;
        PCL_sRegE1      : out    vl_logic;
        PCL_sRegE2      : out    vl_logic;
        PCL_sdqMuxSel   : out    vl_logic;
        PCL_sraRegE1    : out    vl_logic;
        PCL_sraRegE2    : out    vl_logic;
        PCL_srmRegE1    : out    vl_logic;
        PCL_srmRegE2    : out    vl_logic_vector(0 to 2);
        PCL_stSteerCntl : out    vl_logic_vector(0 to 9);
        PCL_timJtgSprHold: out    vl_logic;
        PCL_timSprDcds  : out    vl_logic_vector(0 to 5);
        PCL_tlbRE       : out    vl_logic;
        PCL_tlbSX       : out    vl_logic;
        PCL_tlbWE       : out    vl_logic;
        PCL_tlbWS       : out    vl_logic;
        PCL_trcLoadDV   : out    vl_logic;
        PCL_vctDbgSprHold: out    vl_logic;
        PCL_vctSprDcds  : out    vl_logic_vector(0 to 5);
        PCL_wbAlgnErr   : out    vl_logic;
        PCL_wbClearOrFlush: out    vl_logic;
        PCL_wbClearTerms: out    vl_logic;
        PCL_wbComplete  : out    vl_logic;
        PCL_wbDbgIcmp   : out    vl_logic;
        PCL_wbFullForPO : out    vl_logic;
        PCL_wbFullL2    : out    vl_logic;
        PCL_wbHold      : out    vl_logic;
        PCL_wbHoldNonErr: out    vl_logic;
        PCL_wbLdNotSt   : out    vl_logic;
        PCL_wbRpAddr    : out    vl_logic_vector(0 to 4);
        PCL_wbRpEqdcdApAddr: out    vl_logic;
        PCL_wbRpEqdcdBpAddr: out    vl_logic;
        PCL_wbRpEqdcdSpAddr: out    vl_logic;
        PCL_wbRpWrEn    : out    vl_logic;
        PCL_wbStorageOp : out    vl_logic;
        PCL_wbStrgEnd   : out    vl_logic;
        PCL_xerL2Hold   : out    vl_logic;
        APU_dcdApuOp    : in     vl_logic;
        APU_dcdExeLdDepend: in     vl_logic;
        APU_dcdForceAlgn: in     vl_logic;
        APU_dcdForceBESteering: in     vl_logic;
        APU_dcdFpuOp    : in     vl_logic;
        APU_dcdGprWr    : in     vl_logic;
        APU_dcdLdStByte : in     vl_logic;
        APU_dcdLdStDw   : in     vl_logic;
        APU_dcdLdStHw   : in     vl_logic;
        APU_dcdLdStQw   : in     vl_logic;
        APU_dcdLdStWd   : in     vl_logic;
        APU_dcdLoad     : in     vl_logic;
        APU_dcdLwbLdDepend: in     vl_logic;
        APU_dcdPrivOp   : in     vl_logic;
        APU_dcdRaEn     : in     vl_logic;
        APU_dcdRbEn     : in     vl_logic;
        APU_dcdStore    : in     vl_logic;
        APU_dcdTrapBE   : in     vl_logic;
        APU_dcdTrapLE   : in     vl_logic;
        APU_dcdUpdate   : in     vl_logic;
        APU_dcdWbLdDepend: in     vl_logic;
        APU_dcdXerCAEn  : in     vl_logic;
        APU_dcdXerOVEn  : in     vl_logic;
        APU_exeBlkingMco: in     vl_logic;
        APU_exeBusy     : in     vl_logic;
        APU_exeNonBlkingMco: in     vl_logic;
        CAR_endian      : in     vl_logic;
        CB              : in     vl_logic;
        DBG_dvcRdEn     : in     vl_logic;
        DBG_dvcWrEn     : in     vl_logic;
        DBG_exeIacSuppress: in     vl_logic;
        DBG_icmpEn      : in     vl_logic;
        DBG_wbDacSuppress: in     vl_logic;
        DCU_CA          : in     vl_logic;
        DCU_DA          : in     vl_logic;
        DCU_DOF         : in     vl_logic;
        DCU_carByteEn   : in     vl_logic_vector(0 to 3);
        DCU_firstCycCarStXltV: in     vl_logic;
        DCU_pclOcmLdPendNoWait: in     vl_logic;
        EXE_admMco      : in     vl_logic;
        EXE_divMco      : in     vl_logic;
        EXE_ea          : in     vl_logic_vector(30 to 31);
        EXE_multMco     : in     vl_logic;
        EXE_trap        : in     vl_logic;
        EXE_xerTBC      : in     vl_logic_vector(0 to 6);
        EXE_xerTBCIn    : in     vl_logic_vector(0 to 6);
        EXE_xerTBCNotEqZero: in     vl_logic;
        ICU_LDBE        : in     vl_logic;
        ICU_dsCA        : in     vl_logic;
        ICU_gprDRCC     : in     vl_logic;
        IFB_dcdBubble   : in     vl_logic;
        IFB_dcdDataIn_NEG: in     vl_logic_vector(0 to 31);
        IFB_dcdFull     : in     vl_logic;
        IFB_dcdRegE1    : in     vl_logic;
        IFB_dcdRegE2    : in     vl_logic;
        IFB_exeCorrect  : in     vl_logic;
        IFB_exeFlush    : in     vl_logic;
        IFB_exeRfciL2   : in     vl_logic;
        IFB_exeRfiL2    : in     vl_logic;
        IFB_exeScL2     : in     vl_logic;
        IFB_stepStL2    : in     vl_logic;
        IFB_stuffStL2   : in     vl_logic;
        IFB_trcPipeHold : in     vl_logic;
        LSSD_coreTestEn : in     vl_logic;
        MMU_BMCO        : in     vl_logic;
        MMU_dsStatus    : in     vl_logic_vector(0 to 4);
        MMU_wbHold      : in     vl_logic;
        OCM_DOF         : in     vl_logic;
        OCM_dsComplete  : in     vl_logic;
        PGM_divEn       : in     vl_logic;
        PGM_mmuEn       : in     vl_logic;
        VCT_errorSprSuppress: in     vl_logic;
        VCT_exeSuppForApu: in     vl_logic;
        VCT_exeSuppForCr: in     vl_logic;
        VCT_exeSuppForExe2Clear: in     vl_logic;
        VCT_exeSuppress : in     vl_logic;
        VCT_sxrOR_L2    : in     vl_logic;
        VCT_wbFlush     : in     vl_logic;
        VCT_wbFlushAsync: in     vl_logic;
        VCT_wbLoadSuppress: in     vl_logic;
        VCT_wbSuppress  : in     vl_logic;
        XXX_dcrAck      : in     vl_logic;
        c2Clk           : in     vl_logic;
        coreReset       : in     vl_logic;
        dcdApuValidOp_NEG: in     vl_logic;
        PCL_exeDvcOrParityHold: out    vl_logic;
        ICU_CCR0DPP     : in     vl_logic;
        CAR_cacheable   : in     vl_logic;
        lwbFullL2       : out    vl_logic;
        PCL_lwbCacheableL2: out    vl_logic;
        PCL_dofDregFull : out    vl_logic;
        PCL_BpEqSp      : out    vl_logic;
        PCL_gprRdClk    : out    vl_logic
    );
end p405s_pcl_top;
